.subckt full_bandgap VDD VSS
.ends
.end
