* NGSPICE file created from complete_schematic_pads.ext - technology: ihp-sg13g2

.subckt complete_schematic_pads
X0 a_n7059_10169# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X1 a_981_18638# a_n6059_11418# a_n7415_12373# a_n7415_12373# sg13_lv_nmos ad=0.1005p pd=1.34u as=0.1005p ps=1.34u w=0.15u l=10u
X2 vdd a_n7059_10169# a_n7288_16809# vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X3 a_n7289_16017# a_527_15753# rppd l=38.65u w=0.5u
X4 a_n7288_18340# a_528_18033# rppd l=38.65u w=0.71u
X5 a_n7415_12373# a_5580_15247# a_n7059_10169# a_n7415_12373# sg13_lv_nmos ad=2.448p pd=15.08u as=1.368p ps=7.58u w=7.2u l=9.75u
X6 a_n6059_10861# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X7 a_n7059_10169# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=3.1875p ps=19.43u w=9.375u l=2.08u
X8 a_4707_16560# vdd vdd vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X9 mc_n3216_5326# a_n7415_12373# cap_cmim l=5u w=5u
X10 vdd a_3822_10479# a_n7059_10169# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X11 vdd a_n7059_10169# a_n7288_16809# vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X12 a_6206_12572# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X13 a_5580_15247# a_3630_15211# a_n7415_12373# a_n7415_12373# sg13_lv_nmos ad=0.2448p pd=2.12u as=0.2448p ps=2.12u w=0.72u l=9.75u
X14 vdd a_3822_10479# a_n7059_10169# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X15 vdd a_9247_14192# a_4707_16560# vdd sg13_lv_pmos ad=1.802p pd=11.28u as=1.802p ps=11.28u w=5.3u l=1.95u
X16 a_n7415_12373# a_n6059_10861# a_n6059_11418# a_n7415_12373# sg13_lv_nmos ad=0.33915p pd=2.165u as=0.33915p ps=2.165u w=1.785u l=5u
X17 mc_n7394_8240# a_n7415_12373# cap_cmim l=5u w=5u
X18 a_4238_12572# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=3.1875p ps=19.43u w=9.375u l=2.08u
X19 a_4707_16560# vdd vdd vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X20 vdd a_3822_10479# a_n7059_10169# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X21 vdd a_3822_10479# a_5222_12572# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X22 a_n7288_18340# a_n7415_12373# rppd l=38.65u w=0.71u
X23 vdd a_3822_10479# a_6206_12572# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X24 a_n6059_11418# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X25 mc_n3216_6828# a_n7415_12373# cap_cmim l=5u w=5u
X26 a_n6059_10861# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X27 a_n7415_12373# a_n7289_16545# a_n7289_16545# a_n7415_12373# sg13_lv_nmos ad=0.8925p pd=5.93u as=0.49875p ps=3.005u w=2.625u l=5u
X28 a_1804_15931# a_n7415_12373# cap_cmim l=18.2u w=18.2u
X29 a_n7289_16545# a_n7289_16545# a_n7415_12373# a_n7415_12373# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X30 vdd a_3822_10479# a_4238_12572# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X31 a_n7289_16545# a_n7289_16545# a_n7415_12373# a_n7415_12373# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X32 a_n7289_16017# a_527_16281# rppd l=38.65u w=0.5u
X33 vdd a_n7059_10169# a_n6059_10861# vdd sg13_lv_pmos ad=0.6375p pd=4.43u as=0.35625p ps=2.255u w=1.875u l=5u
X34 a_3630_15211# a_n6059_11418# a_4707_16560# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X35 a_n7059_10169# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X36 a_n6059_11418# a_n6059_10861# a_n7415_12373# a_n7415_12373# sg13_lv_nmos ad=0.33915p pd=2.165u as=0.33915p ps=2.165u w=1.785u l=5u
X37 mc_n4570_8240# a_n7415_12373# cap_cmim l=5u w=5u
X38 a_n7289_16545# a_n7289_16545# a_n7415_12373# a_n7415_12373# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.8925p ps=5.93u w=2.625u l=5u
X39 a_n7288_17727# a_528_18033# rppd l=38.65u w=0.71u
X40 a_n6059_11418# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X41 a_n7288_17115# a_528_16809# rppd l=38.65u w=0.71u
X42 a_n7288_16809# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X43 a_1804_15931# a_981_18638# vdd vdd sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X44 a_5580_15247# a_n6059_10861# a_4707_16560# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X45 a_n7059_10169# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X46 a_n7289_15489# a_527_15753# rppd l=38.65u w=0.5u
X47 a_7190_12572# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X48 vdd a_3822_10479# a_n7059_10169# vdd sg13_lv_pmos ad=3.1875p pd=19.43u as=1.78125p ps=9.755u w=9.375u l=2.08u
X49 vdd a_n7059_10169# a_n6059_11418# vdd sg13_lv_pmos ad=0.6375p pd=4.43u as=0.35625p ps=2.255u w=1.875u l=5u
X50 a_981_18638# a_981_18638# vdd vdd sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X51 a_n7289_15489# a_n6059_10861# rppd l=38.65u w=0.5u
X52 a_n7415_12373# a_n7289_16545# a_n7289_16545# a_n7415_12373# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X53 a_5222_12572# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X54 mc_n1752_8240# a_n7415_12373# cap_cmim l=5u w=5u
X55 mc_n5930_8240# a_n7415_12373# cap_cmim l=5u w=5u
X56 vdd a_3822_10479# a_7190_12572# vdd sg13_lv_pmos ad=3.1875p pd=19.43u as=1.78125p ps=9.755u w=9.375u l=2.08u
X57 a_n7415_12373# a_527_13669# rppd l=38.65u w=3u
X58 a_n7288_16809# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X59 a_n7289_14961# a_n6059_10861# rppd l=38.65u w=0.5u
X60 vdd a_n7059_10169# a_n7288_16809# vdd sg13_lv_pmos ad=0.68p pd=4.68u as=0.38p ps=2.38u w=2u l=5u
X61 a_n6059_11418# a_n6059_10861# a_n7415_12373# a_n7415_12373# sg13_lv_nmos ad=0.33915p pd=2.165u as=0.6069p ps=4.25u w=1.785u l=5u
X62 a_n7415_12373# a_5580_15247# a_n7059_10169# a_n7415_12373# sg13_lv_nmos ad=1.368p pd=7.58u as=1.368p ps=7.58u w=7.2u l=9.75u
X63 a_n6059_10861# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.6375p ps=4.43u w=1.875u l=5u
X64 a_4707_16560# vdd vdd vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X65 mc_n7394_5326# a_n7415_12373# cap_cmim l=5u w=5u
X66 a_n6059_10861# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X67 a_4707_16560# vdd vdd vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X68 mc_n3216_8240# a_n7415_12373# cap_cmim l=5u w=5u
X69 a_n7059_10169# a_5580_15247# a_n7415_12373# a_n7415_12373# sg13_lv_nmos ad=1.368p pd=7.58u as=1.368p ps=7.58u w=7.2u l=9.75u
X70 vdd a_n7059_10169# a_n6059_10861# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X71 a_n6059_11418# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.6375p ps=4.43u w=1.875u l=5u
X72 vdd a_1804_15931# a_n6059_11418# vdd sg13_lv_pmos ad=0.104p pd=1.34u as=0.104p ps=1.34u w=0.2u l=4u
X73 vdd a_981_18638# a_981_18638# vdd sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X74 mc_n7394_6828# a_n7415_12373# cap_cmim l=5u w=5u
X75 a_5580_15247# a_n7059_10169# cap_cmim l=22.29u w=22.29u
X76 a_n6059_11418# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X77 a_5580_15247# a_n6059_10861# a_4707_16560# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X78 vdd a_981_18638# a_1804_15931# vdd sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X79 a_n7415_12373# a_n7289_16545# a_n7289_16545# a_n7415_12373# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X80 a_n7288_17115# a_528_17421# rppd l=38.65u w=0.71u
X81 mc_n4570_5326# a_n7415_12373# cap_cmim l=5u w=5u
X82 a_n7289_16545# a_n7289_16545# a_n7415_12373# a_n7415_12373# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X83 vdd a_n7059_10169# a_n6059_11418# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X84 vdd a_n7059_10169# a_n6059_10861# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X85 a_n7289_14961# a_527_14697# rppd l=38.65u w=0.5u
X86 vdd vdd a_3630_15211# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X87 a_n7415_12373# a_n7289_16545# a_n7289_16545# a_n7415_12373# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X88 a_3630_15211# a_n6059_11418# a_4707_16560# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X89 a_n7288_16809# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.68p ps=4.68u w=2u l=5u
X90 a_n7289_14433# a_527_14697# rppd l=38.65u w=0.5u
X91 vdd a_n7059_10169# a_n6059_10861# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X92 a_n7288_17727# a_528_17421# rppd l=38.65u w=0.71u
X93 mc_n4570_6828# a_n7415_12373# cap_cmim l=5u w=5u
X94 a_n7288_16809# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X95 vdd vdd a_5580_15247# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X96 a_n7288_16809# a_528_16809# rppd l=38.65u w=0.71u
X97 mc_n1752_5326# a_n7415_12373# cap_cmim l=5u w=5u
X98 mc_n5930_5326# a_n7415_12373# cap_cmim l=5u w=5u
X99 a_n7059_10169# a_5580_15247# a_n7415_12373# a_n7415_12373# sg13_lv_nmos ad=1.368p pd=7.58u as=2.448p ps=15.08u w=7.2u l=9.75u
X100 vdd a_n7059_10169# a_n6059_11418# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X101 vdd vdd a_5580_15247# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X102 vdd a_n7059_10169# a_n7288_16809# vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X103 a_n7415_12373# a_n6059_10861# a_n6059_11418# a_n7415_12373# sg13_lv_nmos ad=0.6069p pd=4.25u as=0.33915p ps=2.165u w=1.785u l=5u
X104 a_n7289_16545# a_527_16281# rppd l=38.65u w=0.5u
X105 a_n7289_14433# a_527_13669# rppd l=38.65u w=0.5u
X106 a_3630_15211# a_3630_15211# a_n7415_12373# a_n7415_12373# sg13_lv_nmos ad=0.2448p pd=2.12u as=0.2448p ps=2.12u w=0.72u l=9.75u
X107 vdd a_n7059_10169# a_n6059_11418# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X108 vdd vdd a_3630_15211# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X109 mc_n1752_6828# a_n7415_12373# cap_cmim l=5u w=5u
X110 mc_n5930_6828# a_n7415_12373# cap_cmim l=5u w=5u
C0 a_1804_15931# w_n7489_9836# 0.01614f
C1 vdd w_1450_16710# 0.13483f
C2 mc_n5930_8240# a_n7288_16809# 0.02191f
C3 a_3822_10479# a_n6059_10861# 0.09806f
C4 mc_n5930_6828# mc_n7394_6828# 0.31196f
C5 a_n7203_14433# a_527_13669# 0.01946f
C6 a_n7202_18646# a_n7202_18340# 0.56632f
C7 a_n7059_10169# a_n6059_10861# 3.10863f
C8 vdd mc_n5930_8240# 0.01964f
C9 a_n7203_16017# a_n7289_16017# 0.01946f
C10 a_3630_15211# w_3320_16060# 0.08623f
C11 a_n7289_16545# a_n7202_17727# 0.04493f
C12 mc_n4570_6828# mc_n4570_8240# 0.34633f
C13 a_527_15753# a_n6059_10861# 0.02893f
C14 a_527_16281# a_528_16809# 0.01695f
C15 a_n7203_14961# a_n7289_14961# 0.01946f
C16 mc_n4570_8240# mc_n5930_8240# 0.38921f
C17 a_981_18638# a_n7202_18340# 0.0122f
C18 a_5580_15247# w_3320_10081# 0.01939f
C19 mc_n5930_8240# a_n7059_10169# 0.01546f
C20 a_n7203_15225# a_n7289_14961# 0.01946f
C21 a_n7203_15753# a_n7289_15489# 0.01947f
C22 a_n7203_16017# a_n7289_16545# 0.34937f
C23 a_n7289_16545# a_1804_15931# 0.07823f
C24 a_981_18638# a_n6059_11418# 0.36385f
C25 a_n7203_15753# a_527_15753# 0.01946f
C26 a_527_13669# a_527_14697# 0.01716f
C27 w_1389_15644# a_n6059_11418# 0.01462f
C28 mc_n5930_5326# mc_n5930_6828# 0.29087f
C29 a_n7202_18340# a_n7288_18340# 0.02797f
C30 a_n7203_14433# a_n7203_14697# 0.56632f
C31 vdd w_8745_13831# 0.12219f
C32 a_7190_12572# a_6206_12572# 0.03084f
C33 a_n6059_11418# m3_1900_17599# 0.26018f
C34 a_527_16281# a_527_15753# 0.01716f
C35 mc_n1752_6828# mc_n1752_8240# 0.34633f
C36 a_5580_15247# a_n6059_10861# 1.95475f
C37 a_4707_16560# a_n6059_11418# 1.8134f
C38 vdd a_n7202_18646# 0.09721f
C39 a_n6059_11418# w_n7489_9836# 0.04419f
C40 a_n7289_16545# a_n7289_14961# 0.01076f
C41 w_3320_10081# a_n6059_10861# 0.03529f
C42 vdd a_981_18638# 2.61727f
C43 vdd a_7190_12572# 0.17004f
C44 a_1804_15931# mc_n1752_8240# 0.22161f
C45 vdd a_9247_14192# 1.63687f
C46 vdd w_1389_15644# 0.08151f
C47 a_n7203_14697# a_527_14697# 0.01946f
C48 vdd m3_1900_17599# 0.09884f
C49 vdd a_4707_16560# 3.34935f
C50 w_n7489_9836# a_n7288_16809# 0.03158f
C51 a_7190_12572# a_3822_10479# 4.39984f
C52 a_528_17421# a_n7202_17727# 0.02797f
C53 mc_n5930_8240# mc_n7394_8240# 0.31196f
C54 a_n7289_14433# a_n7289_14961# 0.01716f
C55 vdd w_n7489_9836# 0.42428f
C56 a_1804_15931# mc_n1752_6828# 0.36984f
C57 a_n7289_15489# a_n7203_15489# 0.01947f
C58 mc_n3216_8240# a_n7288_16809# 0.02191f
C59 mc_n4570_6828# mc_n3216_6828# 0.39485f
C60 a_n7289_16545# a_n6059_11418# 0.66075f
C61 a_n7289_16545# a_527_13669# 0.0393f
C62 w_1450_16710# a_n6059_10861# 0.01046f
C63 a_n7288_17727# a_n7288_18340# 0.01705f
C64 a_n7203_14961# a_n7203_14697# 0.56632f
C65 a_n7202_16809# a_n7203_16545# 0.56625f
C66 vdd mc_n3216_8240# 0.01981f
C67 a_n7289_16017# a_n7288_16809# 0.01151f
C68 mc_n3216_5326# mc_n4570_5326# 0.39485f
C69 a_5580_15247# w_8745_13831# 0.01565f
C70 a_6206_12572# a_5222_12572# 0.03081f
C71 mc_n4570_6828# mc_n5930_6828# 0.38921f
C72 w_n7489_9836# a_n7059_10169# 0.0763f
C73 mc_n5930_6828# mc_n5930_8240# 0.34633f
C74 mc_n1752_5326# mc_n3216_5326# 0.31196f
C75 mc_n1752_5326# mc_n1752_6828# 0.29087f
C76 a_n6059_11418# w_3320_16060# 0.0273f
C77 mc_n4570_8240# mc_n3216_8240# 0.39485f
C78 mc_n3216_8240# a_n7059_10169# 0.01528f
C79 a_5222_12572# a_4238_12572# 0.03079f
C80 a_n7289_16545# a_n7288_16809# 0.64582f
C81 a_n6059_11418# a_n7203_13669# 0.02588f
C82 a_n6059_11418# a_3630_15211# 3.28258f
C83 a_n7203_13669# a_527_13669# 0.12082f
C84 vdd a_n7289_16545# 0.36751f
C85 vdd a_5222_12572# 0.16213f
C86 a_n7289_16545# a_n7203_14697# 0.27223f
C87 a_5580_15247# a_9247_14192# 0.0705f
C88 a_n7289_15489# a_n7289_16017# 0.01718f
C89 mc_n1752_5326# a_1804_15931# 0.36984f
C90 a_5580_15247# a_4707_16560# 2.20926f
C91 a_n7202_17115# a_n7289_16545# 0.14683f
C92 a_n7289_16545# a_n7059_10169# 0.19248f
C93 a_3822_10479# a_5222_12572# 4.36409f
C94 vdd w_3320_16060# 0.93176f
C95 a_n7289_15489# a_n7289_16545# 0.01143f
C96 a_528_17421# a_528_18033# 0.01716f
C97 mc_n1752_8240# a_n7288_16809# 0.02191f
C98 vdd a_n7203_13669# 0.01928f
C99 vdd a_3630_15211# 5.84446f
C100 a_n7289_16545# a_527_15753# 0.01192f
C101 vdd mc_n1752_8240# 0.01975f
C102 a_528_17421# a_n6059_11418# 0.01278f
C103 a_n7203_14697# a_n7289_14433# 0.01946f
C104 a_n7203_15489# a_n6059_10861# 0.03922f
C105 a_981_18638# a_n6059_10861# 0.01705f
C106 a_527_14697# a_n6059_10861# 0.0297f
C107 a_n7289_16545# a_n7202_18033# 0.02918f
C108 a_n7203_16017# a_n6059_11418# 0.01623f
C109 w_1389_15644# a_n6059_10861# 0.0227f
C110 a_527_16281# a_n7203_16281# 0.01946f
C111 a_n7289_16545# a_n7202_16809# 0.31907f
C112 a_n6059_11418# a_1804_15931# 1.06328f
C113 a_3630_15211# a_3822_10479# 0.15549f
C114 m3_1900_17599# a_n6059_10861# 0.01692f
C115 w_1450_16710# a_981_18638# 0.01837f
C116 a_527_16281# a_n7203_16545# 0.01946f
C117 a_4707_16560# a_n6059_10861# 1.04184f
C118 a_n7203_15753# a_n7203_15489# 0.56632f
C119 mc_n1752_8240# a_n7059_10169# 0.01528f
C120 vdd mc_n3216_5326# 0.24855f
C121 a_n7289_16545# a_n7202_17421# 0.07627f
C122 w_n7489_9836# a_n6059_10861# 0.01847f
C123 vdd a_n7202_17727# 0.03741f
C124 mc_n3216_6828# mc_n3216_8240# 0.34633f
C125 a_n7203_15225# a_n6059_10861# 0.03934f
C126 a_n7288_17727# a_n7202_17727# 0.02797f
C127 a_528_16809# a_528_17421# 0.01716f
C128 vdd a_1804_15931# 3.95601f
C129 a_n7202_18340# a_528_18033# 0.02797f
C130 a_n7203_16281# a_n7203_16545# 0.56632f
C131 a_5580_15247# w_3320_16060# 0.12191f
C132 vdd mc_n4570_5326# 0.24855f
C133 a_5580_15247# a_3630_15211# 2.48993f
C134 a_n6059_11418# a_528_18033# 0.01068f
C135 w_8745_13831# a_9247_14192# 0.01276f
C136 a_n7289_16545# a_n6059_10861# 0.0901f
C137 a_1804_15931# a_n7059_10169# 0.35354f
C138 a_n7202_18033# a_n7202_17727# 0.56632f
C139 a_981_18638# a_n7202_18646# 0.01155f
C140 vdd mc_n1752_5326# 0.24855f
C141 a_3630_15211# w_3320_10081# 0.01456f
C142 a_n6059_11418# a_527_13669# 0.01087f
C143 vdd mc_n7394_5326# 0.47046f
C144 a_4707_16560# w_8745_13831# 0.01171f
C145 a_n7203_16017# a_527_15753# 0.01946f
C146 mc_n7394_5326# mc_n7394_6828# 0.29087f
C147 a_n7203_15753# a_n7289_16545# 0.3003f
C148 a_n7202_18646# a_n7288_18340# 0.02797f
C149 w_3320_16060# a_n6059_10861# 0.06145f
C150 a_n7202_17421# a_n7202_17727# 0.56632f
C151 a_527_16281# a_n7289_16545# 0.03573f
C152 a_n7289_15489# a_n7289_14961# 0.01718f
C153 a_3630_15211# a_n6059_10861# 2.21895f
C154 vdd a_n7202_18340# 0.0576f
C155 a_528_17421# a_n7202_17421# 0.02797f
C156 a_981_18638# m3_1900_17599# 0.06332f
C157 mc_n5930_5326# mc_n4570_5326# 0.38921f
C158 a_4707_16560# a_9247_14192# 0.52791f
C159 vdd a_n6059_11418# 6.78922f
C160 a_n7289_16017# a_n7203_16281# 0.01946f
C161 a_5580_15247# a_1804_15931# 1.05678f
C162 a_n7203_14961# a_527_14697# 0.01946f
C163 a_n7203_15225# a_n7203_15489# 0.56632f
C164 a_528_16809# a_n6059_11418# 0.02012f
C165 vdd a_6206_12572# 0.16195f
C166 a_n7289_16545# a_n7203_14433# 0.28328f
C167 mc_n5930_5326# mc_n7394_5326# 0.31196f
C168 mc_n3216_5326# mc_n3216_6828# 0.29087f
C169 mc_n1752_6828# mc_n3216_6828# 0.31196f
C170 a_n6059_11418# a_n7059_10169# 2.78705f
C171 a_n7289_16545# a_n7203_16281# 0.46335f
C172 vdd a_4238_12572# 0.16979f
C173 a_3822_10479# a_6206_12572# 4.40911f
C174 a_n7289_16545# a_n7203_16545# 0.57323f
C175 vdd a_n7288_16809# 2.7233f
C176 a_n7202_18340# a_n7202_18033# 0.5628f
C177 a_n7202_18033# a_528_18033# 0.02797f
C178 a_n7288_17115# a_n7288_16809# 0.0308f
C179 a_n6059_11418# a_527_15753# 0.01738f
C180 a_n7203_14961# a_n7203_15225# 0.56632f
C181 a_1804_15931# a_n6059_10861# 0.63328f
C182 a_n7289_16545# a_n7203_15489# 0.27748f
C183 a_3822_10479# a_4238_12572# 4.39975f
C184 a_n7203_14433# a_n7203_13669# 0.56632f
C185 a_n7289_16545# a_527_14697# 0.01226f
C186 vdd mc_n7394_6828# 0.22191f
C187 a_n7203_14433# a_n7289_14433# 0.01946f
C188 mc_n4570_8240# a_n7288_16809# 0.02191f
C189 a_n7059_10169# a_n7288_16809# 10.5491f
C190 a_n7202_16809# a_n6059_11418# 0.03367f
C191 a_n7203_15753# a_n7203_16017# 0.56632f
C192 w_1450_16710# a_1804_15931# 0.02886f
C193 vdd a_3822_10479# 51.183f
C194 a_n7288_17727# a_n7288_17115# 0.01716f
C195 vdd mc_n4570_8240# 0.01975f
C196 a_n7289_15489# a_n7288_16809# 0.01126f
C197 vdd a_n7059_10169# 53.0636f
C198 a_n7202_17115# a_n7288_17115# 0.02797f
C199 a_n7202_17115# a_528_16809# 0.02797f
C200 a_n6059_11418# a_n7202_17421# 0.01101f
C201 a_5580_15247# a_n6059_11418# 0.66736f
C202 a_n7289_16545# w_n7489_9836# 0.04233f
C203 mc_n4570_6828# mc_n4570_5326# 0.29087f
C204 a_n7289_16545# a_n7203_14961# 0.25927f
C205 vdd a_527_15753# 0.01523f
C206 a_n7289_16545# a_n7203_15225# 0.26585f
C207 a_3822_10479# a_n7059_10169# 3.82737f
C208 mc_n4570_8240# a_n7059_10169# 0.01528f
C209 a_n7202_16809# a_n7288_16809# 0.06913f
C210 vdd a_n7202_18033# 0.04632f
C211 vdd mc_n5930_5326# 0.24855f
C212 a_4707_16560# w_3320_16060# 0.05243f
C213 a_n7289_16545# a_n7289_16017# 0.03605f
C214 a_4707_16560# a_3630_15211# 2.47471f
C215 a_528_16809# a_n7202_16809# 0.02797f
C216 a_n7288_17727# a_n7202_18033# 0.02797f
C217 a_n7203_16017# a_n7203_16281# 0.56632f
C218 vdd a_5580_15247# 10.1146f
C219 a_n7202_17115# a_n7202_16809# 0.56632f
C220 a_n7288_17115# a_n7202_17421# 0.02797f
C221 a_n6059_11418# a_n6059_10861# 8.04164f
C222 mc_n7394_8240# a_n7288_16809# 0.02191f
C223 vdd w_3320_10081# 0.29549f
C224 mc_n1752_8240# mc_n3216_8240# 0.31196f
C225 w_1450_16710# a_n6059_11418# 0.02162f
C226 a_n7202_17115# a_n7202_17421# 0.56632f
C227 a_5580_15247# a_3822_10479# 0.02769f
C228 vdd mc_n7394_8240# 0.24657f
C229 a_5580_15247# a_n7059_10169# 32.0404f
C230 a_4238_12572# a_n6059_10861# 0.01263f
C231 a_981_18638# a_1804_15931# 1.49127f
C232 mc_n7394_6828# mc_n7394_8240# 0.34633f
C233 w_1389_15644# a_1804_15931# 0.04245f
C234 w_3320_10081# a_3822_10479# 0.03683f
C235 a_n6059_10861# a_n7288_16809# 1.54398f
C236 w_3320_10081# a_n7059_10169# 0.03712f
C237 a_n7289_16545# a_n7203_13669# 2.15576f
C238 a_1804_15931# m3_1900_17599# 0.19321f
C239 vdd a_n6059_10861# 7.9717f
C240 a_n7289_16545# a_n7289_14433# 0.01035f
C241 mc_n7394_8240# a_n7059_10169# 0.01052f
C242 mc_n1752_5326# a_n7415_12373# 1.92145f $ **FLOATING
C243 mc_n3216_5326# a_n7415_12373# 1.85536f $ **FLOATING
C244 mc_n4570_5326# a_n7415_12373# 1.86279f $ **FLOATING
C245 mc_n5930_5326# a_n7415_12373# 1.85511f $ **FLOATING
C246 mc_n7394_5326# a_n7415_12373# 1.86582f $ **FLOATING
C247 mc_n1752_6828# a_n7415_12373# 1.89719f $ **FLOATING
C248 mc_n3216_6828# a_n7415_12373# 1.83111f $ **FLOATING
C249 mc_n4570_6828# a_n7415_12373# 1.83853f $ **FLOATING
C250 mc_n5930_6828# a_n7415_12373# 1.83085f $ **FLOATING
C251 mc_n7394_6828# a_n7415_12373# 1.84156f $ **FLOATING
C252 mc_n1752_8240# a_n7415_12373# 2.05251f $ **FLOATING
C253 mc_n3216_8240# a_n7415_12373# 1.93901f $ **FLOATING
C254 mc_n4570_8240# a_n7415_12373# 1.94644f $ **FLOATING
C255 mc_n5930_8240# a_n7415_12373# 1.93875f $ **FLOATING
C256 mc_n7394_8240# a_n7415_12373# 1.94947f $ **FLOATING
C257 m3_1900_17599# a_n7415_12373# 0.07285f
C258 a_7190_12572# a_n7415_12373# 0.15504f $ **FLOATING
C259 a_6206_12572# a_n7415_12373# 0.10855f $ **FLOATING
C260 a_5222_12572# a_n7415_12373# 0.10229f $ **FLOATING
C261 a_4238_12572# a_n7415_12373# 0.13225f $ **FLOATING
C262 a_3822_10479# a_n7415_12373# 13.9081f $ **FLOATING
C263 a_n7059_10169# a_n7415_12373# 18.8682f $ **FLOATING
C264 a_n7203_13669# a_n7415_12373# 13.2663f
C265 a_527_13669# a_n7415_12373# 0.57989f $ **FLOATING
C266 a_n7203_14433# a_n7415_12373# 3.81224f
C267 a_n7203_14697# a_n7415_12373# 3.80746f
C268 a_n7289_14433# a_n7415_12373# 0.26883f $ **FLOATING
C269 a_9247_14192# a_n7415_12373# 0.87526f $ **FLOATING
C270 a_527_14697# a_n7415_12373# 0.25188f $ **FLOATING
C271 a_n7203_14961# a_n7415_12373# 3.80233f
C272 a_n7203_15225# a_n7415_12373# 3.79878f
C273 a_n7289_14961# a_n7415_12373# 0.25151f $ **FLOATING
C274 a_n7203_15489# a_n7415_12373# 3.79878f
C275 a_n7203_15753# a_n7415_12373# 3.79878f
C276 a_n7289_15489# a_n7415_12373# 0.25183f $ **FLOATING
C277 a_527_15753# a_n7415_12373# 0.23297f $ **FLOATING
C278 a_n7203_16017# a_n7415_12373# 3.79878f
C279 a_n7203_16281# a_n7415_12373# 3.79878f
C280 a_n7289_16017# a_n7415_12373# 0.25124f $ **FLOATING
C281 a_3630_15211# a_n7415_12373# 6.36779f $ **FLOATING
C282 a_5580_15247# a_n7415_12373# 51.7544f $ **FLOATING
C283 a_4707_16560# a_n7415_12373# 1.69969f $ **FLOATING
C284 a_n6059_10861# a_n7415_12373# 15.1337f $ **FLOATING
C285 a_1804_15931# a_n7415_12373# 20.0144f $ **FLOATING
C286 a_n6059_11418# a_n7415_12373# 9.66571f $ **FLOATING
C287 a_527_16281# a_n7415_12373# 0.28604f $ **FLOATING
C288 a_n7203_16545# a_n7415_12373# 3.79788f
C289 a_n7289_16545# a_n7415_12373# 36.4829f $ **FLOATING
C290 a_n7202_16809# a_n7415_12373# 4.50753f
C291 a_n7288_16809# a_n7415_12373# 3.39149f $ **FLOATING
C292 a_528_16809# a_n7415_12373# 0.34584f $ **FLOATING
C293 a_n7202_17115# a_n7415_12373# 4.50921f
C294 a_n7202_17421# a_n7415_12373# 4.50921f
C295 a_n7288_17115# a_n7415_12373# 0.30345f $ **FLOATING
C296 a_528_17421# a_n7415_12373# 0.34565f $ **FLOATING
C297 a_n7202_17727# a_n7415_12373# 4.50921f
C298 a_n7202_18033# a_n7415_12373# 4.51745f
C299 a_n7288_17727# a_n7415_12373# 0.30438f $ **FLOATING
C300 a_528_18033# a_n7415_12373# 0.36381f $ **FLOATING
C301 a_n7202_18340# a_n7415_12373# 4.55105f
C302 a_981_18638# a_n7415_12373# 1.17046f $ **FLOATING
C303 a_n7202_18646# a_n7415_12373# 5.27974f
C304 a_n7288_18340# a_n7415_12373# 0.3202f $ **FLOATING
C305 w_n7489_9836# a_n7415_12373# 0.21456f
C306 w_3320_10081# a_n7415_12373# 0.1031f
C307 w_8745_13831# a_n7415_12373# 0.02418f
C308 w_3320_16060# a_n7415_12373# 0.123f
C309 w_1450_16710# a_n7415_12373# 0.03111f
C310 vdd a_n7415_12373# 69.7956f $ **FLOATING
.ends
