** sch_path: /foss/designs/thesis/thesis_hp/designs/otas/1_schematics/foldedcascode_nmos.sch
.subckt foldedcascode_nmos AVDD PLUS MINUS Vout Ibias d_ena AVSS
*.PININFO AVSS:I Ibias:I AVDD:I PLUS:I MINUS:I Vout:O d_ena:I
XMb net16 net1 AVSS AVSS sg13_lv_nmos w=5u l=5u ng=1 m=1
XMpd5 net1 ena_n AVSS AVSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMpd6 net16 ena net1 AVSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMb1 net14 net1 AVSS AVSS sg13_lv_nmos w=5u l=5u ng=1 m=1
Vmeas net15 net14 0
.save i(vmeas)
XM11 net15 net3 net2 AVDD sg13_lv_pmos w=11.5u l=1.5u ng=2 m=1
XM12 net2 net2 AVDD AVDD sg13_lv_pmos w=11.5u l=1.5u ng=2 m=1
XM18 AVSS net3 net6 AVDD sg13_lv_pmos w=15u l=0.5u ng=5 m=1
XM17 net6 net2 AVDD AVDD sg13_lv_pmos w=11.5u l=1.5u ng=2 m=1
XM9 net5 net2 AVDD AVDD sg13_lv_pmos w=11.5u l=1.5u ng=2 m=1
XM5 net3 net6 net5 AVDD sg13_lv_pmos w=11u l=1.5u ng=2 m=1
XM7 net3 net13 net4 AVSS sg13_lv_nmos w=3u l=2u ng=1 m=1
XM3 net4 net3 AVSS AVSS sg13_lv_nmos w=2.5u l=2u ng=1 m=1
XMpd7 net2 ena AVDD AVDD sg13_lv_pmos w=1u l=0.13u ng=1 m=1
XMpd8 net6 ena AVDD AVDD sg13_lv_pmos w=1u l=0.13u ng=1 m=1
XMt net7 net1 AVSS AVSS sg13_lv_nmos w=5u l=5u ng=1 m=1
XM1 net5 PLUS net7 AVSS sg13_lv_nmos w=6u l=1u ng=1 m=1
XM2 net8 MINUS net7 AVSS sg13_lv_nmos w=6u l=1u ng=1 m=1
XM6 Vout net6 net8 AVDD sg13_lv_pmos w=11u l=1.5u ng=2 m=1
XM0 net8 net2 AVDD AVDD sg13_lv_pmos w=11.5u l=1.5u ng=2 m=1
XMdecoup3 AVDD net2 AVDD AVDD sg13_lv_pmos w=12u l=0.5u ng=4 m=1
XMdecoup4 AVDD net6 AVDD AVDD sg13_lv_pmos w=12u l=0.5u ng=4 m=1
XM8 Vout net13 net9 AVSS sg13_lv_nmos w=3u l=2u ng=1 m=1
XM4 net9 net3 AVSS AVSS sg13_lv_nmos w=2.5u l=2u ng=1 m=1
XMdecoup1 AVSS net1 AVSS AVSS sg13_lv_nmos w=8u l=1u ng=4 m=1
XM13 net10 net2 AVDD AVDD sg13_lv_pmos w=11.5u l=1.5u ng=2 m=1
Vmeas2 net10 net11 0
.save i(vmeas2)
XM15 net11 Vout net12 AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
XM16 net12 net12 AVSS AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
XM14 net13 net12 AVSS AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
XM10 AVDD Vout net13 AVSS sg13_lv_nmos w=15u l=0.5u ng=5 m=1
XMpd11 Vout ena_n AVSS AVSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMdecoup2 AVSS net13 AVSS AVSS sg13_lv_nmos w=8u l=1u ng=4 m=1
XMpd10 net13 ena_n AVSS AVSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMpd9 net3 ena_n AVSS AVSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMpd2 ena_n d_ena AVDD AVDD sg13_lv_pmos w=1u l=0.13u ng=1 m=1
Vmeas1 Ibias net16 0
.save i(vmeas1)
XMpd3 ena ena_n AVDD AVDD sg13_lv_pmos w=1u l=0.13u ng=1 m=1
XMpd1 ena_n d_ena AVSS AVSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XMpd4 ena ena_n AVSS AVSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
.ends
