.subckt complete_schematic_pads_fillers VDD VSS
.ends
.end
