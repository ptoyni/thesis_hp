* Extracted by KLayout with SG13G2 LVS runset on : 16/07/2025 02:34

.SUBCKT ota_final AVSS PLUS AVDD VOUT IBIAS MINUS
M$1 AVDD VOUT \$18643 AVSS sg13_lv_nmos L=0.5u W=15u AS=3.4125p AD=3.4125p
+ PS=20.57u PD=20.57u
M$5 AVSS IBIAS IBIAS AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$9 AVSS IBIAS \$19588 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$13 AVSS IBIAS \$19587 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$17 AVSS AVSS \$19749 AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$18 \$19749 MINUS \$19587 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p
+ PS=6.76u PD=6.76u
M$19 \$19587 PLUS \$19750 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p
+ PS=6.76u PD=6.76u
M$20 \$19750 AVSS AVSS AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$25 \$19588 \$19202 \$19694 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
M$29 AVSS \$19202 \$19695 AVDD sg13_lv_pmos L=0.5u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
C$33 VOUT AVSS cap_cmim w=25.82u l=25.82u A=666.6724p P=103.28u m=1
M$34 \$18645 VOUT \$18646 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$36 AVSS AVSS \$18645 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$37 \$18645 \$18645 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$38 AVSS \$18645 \$18643 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$42 AVDD AVDD \$19694 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p
+ PS=11.56u PD=11.56u
M$43 \$19694 \$19694 AVDD AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$44 AVDD \$19694 \$19695 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$46 AVDD \$19694 \$18646 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$56 AVSS AVSS VOUT AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$57 VOUT \$18643 \$I485994 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$60 AVSS AVSS \$I485993 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$61 \$I485993 \$19202 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$64 AVSS AVSS \$I485994 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$65 \$I485994 \$19202 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$68 AVSS AVSS \$19202 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$69 \$19202 \$18643 \$I485993 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$72 AVDD AVDD \$19202 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p
+ PS=11.56u PD=11.56u
M$73 \$19202 \$19695 \$19750 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$78 AVDD AVDD VOUT AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$79 VOUT \$19695 \$19749 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$84 AVDD AVDD \$19749 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
M$86 AVDD \$19694 \$19750 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$88 AVDD \$19694 \$19749 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
.ENDS ota_final
