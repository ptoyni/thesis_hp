* NGSPICE file created from foldedcascode_nmos_withdummies.ext - technology: ihp-sg13g2

.subckt foldedcascode_nmos_withdummies PLUS MINUS VOUT AVSS AVDD IBIAS D_ENA
X0 AVSS AVSS a_n686_n3376# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X1 AVSS a_n13165_n3086# AVSS AVSS sg13_lv_nmos ad=0.38p pd=2.38u as=0.2167n ps=1.39985m w=2u l=1u
X2 AVDD a_n2227_3805# AVDD AVDD sg13_lv_pmos ad=1.02p pd=6.68u as=0.19842n ps=1.23365m w=3u l=1u
X3 a_492_n6342# AVSS AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X4 AVSS a_n13165_n3086# a_n9134_n1298# AVSS sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X5 a_n13597_n4844# D_ENA AVDD AVDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=0.13u
X6 a_7669_2986# a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X7 AVSS AVSS a_n686_n5390# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X8 a_n2559_1528# a_n8239_n7963# a_n9134_n2395# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X9 a_7669_5842# a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X10 AVDD a_n2559_1528# a_n2343_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X11 a_n722_n4252# VOUT AVDD AVSS sg13_lv_nmos ad=0.7125p pd=4.13u as=1.275p ps=8.18u w=3.75u l=0.5u
X12 AVSS a_n722_n4252# AVSS AVSS sg13_lv_nmos ad=0.68p pd=4.68u as=0 ps=0 w=2u l=1u
X13 AVDD a_n2559_1528# a_n2343_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X14 AVSS AVSS a_n2343_7081# AVSS sg13_lv_nmos ad=1.02p pd=6.68u as=0.57p ps=3.38u w=3u l=1u
X15 AVDD a_n2835_1528# AVDD AVDD sg13_lv_pmos ad=1.02p pd=6.68u as=0 ps=0 w=3u l=1u
X16 a_n722_n4252# VOUT AVDD AVSS sg13_lv_nmos ad=0.7125p pd=4.13u as=0.7125p ps=4.13u w=3.75u l=0.5u
X17 a_7578_n5569# AVSS AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X18 a_7669_1082# AVDD AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X19 a_n686_n6342# AVSS AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X20 AVSS AVSS a_n1391_7081# AVSS sg13_lv_nmos ad=1.02p pd=6.68u as=0.57p ps=3.38u w=3u l=1u
X21 AVSS a_n8239_n7963# a_n2227_3805# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=0.5u
X22 a_7669_3938# a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X23 IBIAS a_n13165_n3086# AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X24 a_1623_5158# a_n2227_3805# a_1623_4682# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X25 AVDD AVDD a_7669_6794# AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X26 AVSS AVSS a_7578_n5569# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X27 AVSS a_n13165_n3086# IBIAS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X28 AVDD a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=1u
X29 a_n2191_4681# a_n2227_3805# a_n2191_4205# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X30 a_n9134_n1298# a_n13165_n3086# AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X31 a_n2191_4205# a_n2227_3805# a_n8239_n7963# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X32 AVSS a_n722_n4252# AVSS AVSS sg13_lv_nmos ad=0.38p pd=2.38u as=0 ps=0 w=2u l=1u
X33 a_n2343_7081# a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X34 AVDD AVDD a_n2343_7081# AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X35 a_n2343_7081# AVDD AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X36 a_n13561_n4818# a_n13597_n4844# AVSS AVSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=0.13u
X37 AVSS a_n13165_n3086# IBIAS AVSS sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X38 a_n9134_n2395# a_n8239_n7963# a_n2559_1528# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X39 a_492_n5866# a_n8239_n7963# a_492_n6342# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X40 a_n8239_n7963# a_n13597_n4844# AVSS AVSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=0.13u
X41 a_492_n3852# a_n722_n4252# a_492_n4328# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X42 AVDD a_n2559_1528# a_7669_4890# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X43 AVDD a_n2559_1528# a_n1391_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X44 AVDD a_n2559_1528# a_7669_2034# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X45 VOUT AVDD AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X46 a_n1391_7081# a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X47 AVSS a_7578_n5569# a_7578_n5569# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X48 a_n2559_1528# a_n8239_n7963# a_n9134_n2395# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X49 a_n1391_7081# AVSS AVSS AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=1.02p ps=6.68u w=3u l=1u
X50 a_n8239_n7963# a_n2227_3805# a_n2191_5157# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X51 a_n2227_3805# a_n8239_n7963# AVSS AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=0.5u
X52 a_n686_n5866# a_n8239_n7963# a_n686_n6342# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X53 AVSS a_n8239_n7963# a_n2227_3805# AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=0.5u
X54 AVDD a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=1u
X55 a_n686_n3852# a_n722_n4252# a_n686_n4328# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X56 a_7578_n5569# VOUT a_9374_n4648# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X57 a_n13165_n3086# a_n13561_n4818# IBIAS AVSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=0.13u
X58 AVDD a_n2227_3805# AVDD AVDD sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=1u
X59 a_8530_n5569# a_7578_n5569# AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X60 AVSS a_n13165_n3086# AVSS AVSS sg13_lv_nmos ad=0.38p pd=2.38u as=0 ps=0 w=2u l=1u
X61 a_n9134_n1298# MINUS a_n1391_7081# AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X62 AVDD a_n2559_1528# a_7669_5842# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X63 a_7669_6794# a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X64 IBIAS a_n13165_n3086# AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X65 a_492_n5390# a_n8239_n7963# a_492_n5866# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X66 AVSS a_n722_n4252# AVSS AVSS sg13_lv_nmos ad=0.38p pd=2.38u as=0 ps=0 w=2u l=1u
X67 a_n9134_n2395# a_n8239_n7963# a_n2559_1528# AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X68 a_n8239_n7963# AVDD AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X69 a_492_n3376# a_n722_n4252# a_492_n3852# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X70 AVDD VOUT a_n722_n4252# AVSS sg13_lv_nmos ad=1.275p pd=8.18u as=0.7125p ps=4.13u w=3.75u l=0.5u
X71 a_n9134_n2395# a_n13165_n3086# AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X72 AVSS a_n13165_n3086# AVSS AVSS sg13_lv_nmos ad=0.38p pd=2.38u as=0 ps=0 w=2u l=1u
X73 AVSS a_n13165_n3086# a_n9134_n2395# AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X74 a_n2343_7081# PLUS a_n9134_n1298# AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X75 a_7669_2034# a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X76 AVDD a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=1u
X77 a_n2343_7081# AVDD AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X78 AVSS a_n2937_n2952# AVSS AVSS sg13_lv_nmos ad=0.68p pd=4.68u as=0 ps=0 w=2u l=1u
X79 AVSS a_n13165_n3086# a_n9134_n2395# AVSS sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X80 a_n2191_5157# a_n2227_3805# a_n2191_4681# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X81 AVDD AVDD VOUT AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X82 a_n686_n5390# a_n8239_n7963# a_n686_n5866# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X83 a_n13597_n4844# D_ENA AVSS AVSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=0.13u
X84 a_n2227_3805# a_n8239_n7963# AVSS AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=0.5u
X85 a_n686_n3376# a_n722_n4252# a_n686_n3852# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X86 a_n2343_7081# a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X87 AVDD a_n2559_1528# a_n1391_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X88 a_492_n4328# AVSS AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X89 a_7578_n5569# a_7578_n5569# AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X90 AVDD VOUT a_n722_n4252# AVSS sg13_lv_nmos ad=0.7125p pd=4.13u as=0.7125p ps=4.13u w=3.75u l=0.5u
X91 AVDD a_n2559_1528# a_7669_2986# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X92 a_1623_4206# a_n2227_3805# VOUT AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X93 a_1623_4682# a_n2227_3805# a_1623_4206# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X94 AVDD AVDD a_n8239_n7963# AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X95 AVSS AVSS a_492_n3376# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X96 a_n2343_7081# AVSS AVSS AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=1.02p ps=6.68u w=3u l=1u
X97 AVDD a_n2227_3805# AVDD AVDD sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=1u
X98 AVDD AVDD a_n2343_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X99 AVSS AVSS a_492_n5390# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X100 a_n9134_n2395# a_n13165_n3086# AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X101 a_n686_n4328# AVSS AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X102 AVDD a_n2559_1528# a_7669_1082# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X103 a_n13561_n4818# a_n13597_n4844# AVDD AVDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=0.13u
X104 a_7669_4890# a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X105 a_n9134_n1298# a_n13165_n3086# AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X106 a_n1391_7081# a_n2559_1528# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X107 a_9374_n4648# VOUT a_7578_n5569# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X108 AVSS a_n722_n4252# AVSS AVSS sg13_lv_nmos ad=0.38p pd=2.38u as=0 ps=0 w=2u l=1u
X109 a_n1391_7081# MINUS a_n9134_n1298# AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X110 AVSS a_n13165_n3086# a_n9134_n1298# AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X111 a_n9134_n1298# PLUS a_n2343_7081# AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X112 AVDD a_n2227_3805# AVDD AVDD sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=1u
X113 AVDD a_n2559_1528# a_7669_3938# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X114 VOUT a_n2227_3805# a_1623_5158# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X115 AVSS a_7578_n5569# a_8530_n5569# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
C0 a_n8239_n7963# a_n722_n4252# 0.50656f
C1 a_n686_n5390# m1_n686_n6334# 0.03177f
C2 VOUT a_n8239_n7963# 0.24186f
C3 VOUT a_n722_n4252# 1.13562f
C4 a_n2559_1528# a_n1391_7081# 0.97281f
C5 a_n2343_7081# a_1623_4206# 0.07239f
C6 a_n2559_1528# a_n2343_7081# 1.444f
C7 a_n2559_1528# a_n2835_1528# 0.062f
C8 a_n13597_n4844# IBIAS 0.10477f
C9 a_n9134_n1298# a_n9134_n2395# 0.0392f
C10 a_n13165_n3086# AVDD 0.01192f
C11 a_n1391_7081# a_n8239_n7963# 0.24946f
C12 a_n2227_3805# AVDD 15.5067f
C13 a_n2343_7081# VOUT 0.2467f
C14 a_n2343_7081# a_1623_5158# 0.07216f
C15 a_n9134_n2395# a_n13165_n3086# 1.3416f
C16 a_n13561_n4818# IBIAS 0.08911f
C17 D_ENA AVDD 0.30593f
C18 a_9374_n4648# a_n2227_3805# 0.10225f
C19 a_n9134_n2395# a_n2227_3805# 0.11372f
C20 a_n686_n3376# a_n8239_n7963# 0.03238f
C21 a_8530_n5569# a_n722_n4252# 0.03137f
C22 PLUS a_n1391_7081# 0.35705f
C23 a_n2343_7081# PLUS 0.31437f
C24 m1_492_n6334# a_492_n3852# 0.03122f
C25 a_n2343_7081# a_n1391_7081# 0.36088f
C26 a_9374_n4648# a_7669_2986# 0.06823f
C27 a_7669_2034# a_n2227_3805# 0.07179f
C28 a_n9134_n1298# a_n8239_n7963# 0.09814f
C29 m1_492_n6334# a_492_n5390# 0.03183f
C30 a_9374_n4648# AVDD 1.21514f
C31 a_n9134_n2395# AVDD 2.31589f
C32 a_n2559_1528# a_7669_1082# 0.0746f
C33 a_n2559_1528# a_n2227_3805# 1.26946f
C34 a_n686_n6342# m1_n686_n6334# 0.03135f
C35 a_n1391_7081# a_n2191_4205# 0.07238f
C36 a_n2559_1528# a_7669_6794# 0.06988f
C37 a_n13165_n3086# a_n8239_n7963# 0.16456f
C38 D_ENA a_n13597_n4844# 0.18618f
C39 a_n9134_n1298# PLUS 0.23501f
C40 a_n9134_n1298# a_n1391_7081# 0.1784f
C41 a_n13561_n4818# a_n13165_n3086# 0.0201f
C42 a_n13597_n4844# AVDD 0.68317f
C43 a_n2227_3805# a_n8239_n7963# 1.43165f
C44 a_n2343_7081# a_n9134_n1298# 0.23934f
C45 a_7669_5842# a_n2227_3805# 0.06914f
C46 a_n2559_1528# AVDD 29.6208f
C47 VOUT a_492_n3376# 0.03213f
C48 VOUT a_n2227_3805# 1.19253f
C49 MINUS PLUS 0.25746f
C50 MINUS a_n1391_7081# 0.51932f
C51 a_n2343_7081# MINUS 0.23141f
C52 a_n8239_n7963# AVDD 7.10925f
C53 a_9374_n4648# a_n2559_1528# 0.83984f
C54 AVDD a_n722_n4252# 0.91757f
C55 a_n2559_1528# a_n9134_n2395# 0.32102f
C56 a_n13561_n4818# AVDD 0.39016f
C57 VOUT AVDD 2.66834f
C58 a_n686_n4328# a_n8239_n7963# 0.03197f
C59 a_n1391_7081# a_n2227_3805# 1.01797f
C60 a_9374_n4648# a_7578_n5569# 0.11814f
C61 a_n2343_7081# a_n2227_3805# 1.18866f
C62 a_n13165_n3086# IBIAS 1.0955f
C63 a_9374_n4648# a_n8239_n7963# 0.01919f
C64 a_n9134_n2395# a_n8239_n7963# 1.17252f
C65 a_9374_n4648# VOUT 0.26312f
C66 m1_n686_n6334# a_n8239_n7963# 0.4315f
C67 VOUT a_n9134_n2395# 0.20229f
C68 m1_492_n6334# a_492_n6342# 0.03137f
C69 m1_n686_n6334# a_n722_n4252# 0.23704f
C70 MINUS a_n9134_n1298# 0.25143f
C71 a_n1391_7081# AVDD 2.24503f
C72 a_n2937_n2952# a_n13165_n3086# 0.07791f
C73 a_9374_n4648# a_7669_4890# 0.06998f
C74 a_n2343_7081# AVDD 3.61544f
C75 a_n2835_1528# AVDD 0.65631f
C76 VOUT a_1623_4682# 0.07308f
C77 IBIAS AVDD 0.16629f
C78 a_n9134_n1298# a_n13165_n3086# 1.52604f
C79 a_n2559_1528# a_7669_3938# 0.07097f
C80 a_n13597_n4844# a_n8239_n7963# 0.05059f
C81 a_492_n4328# VOUT 0.03151f
C82 a_n9134_n2395# a_n1391_7081# 0.06215f
C83 a_n13561_n4818# a_n13597_n4844# 0.1902f
C84 a_n2559_1528# a_n8239_n7963# 1.01131f
C85 a_n2343_7081# a_n9134_n2395# 0.06236f
C86 a_n1391_7081# a_n2191_5157# 0.07207f
C87 m1_492_n6334# a_n8239_n7963# 0.28698f
C88 a_n8239_n7963# a_n2191_4681# 0.07259f
C89 m1_492_n6334# a_n722_n4252# 0.30261f
C90 m1_492_n6334# VOUT 0.10634f
C91 a_7578_n5569# a_n722_n4252# 0.27985f
C92 a_n686_n3852# m1_n686_n6334# 0.03124f
C93 VOUT a_7578_n5569# 0.33361f
C94 D_ENA AVSS 6.65333f
C95 IBIAS AVSS 8.87644f
C96 PLUS AVSS 3.30848f
C97 MINUS AVSS 2.83276f
C98 VOUT AVSS 16.5276f
C99 AVDD AVSS 40.6103f
C100 m1_492_n6334# AVSS 1.43209f
C101 m1_n686_n6334# AVSS 1.40245f
C102 a_492_n5866# AVSS 0.03034f $ **FLOATING
C103 a_n686_n5866# AVSS 0.03052f $ **FLOATING
C104 a_9374_n4648# AVSS 4.05743f $ **FLOATING
C105 a_7578_n5569# AVSS 4.70064f $ **FLOATING
C106 a_n13597_n4844# AVSS 4.03323f $ **FLOATING
C107 a_n2937_n2952# AVSS 0.70555f $ **FLOATING
C108 a_n722_n4252# AVSS 11.4468f $ **FLOATING
C109 a_n13561_n4818# AVSS 1.56383f $ **FLOATING
C110 a_n9134_n2395# AVSS 6.75069f $ **FLOATING
C111 a_n13165_n3086# AVSS 32.2105f $ **FLOATING
C112 a_n9134_n1298# AVSS 3.32115f $ **FLOATING
C113 a_n2835_1528# AVSS 0.28088f $ **FLOATING
C114 a_n2227_3805# AVSS 8.85767f $ **FLOATING
C115 a_n8239_n7963# AVSS 19.7524f $ **FLOATING
C116 a_n1391_7081# AVSS 3.87171f $ **FLOATING
C117 a_n2343_7081# AVSS 2.29815f $ **FLOATING
C118 a_n2559_1528# AVSS 14.1048f $ **FLOATING
.ends
