** sch_path: /foss/designs/thesis_hp/designs/otas/1_schematics/foldedcascode_nmos_withdummies.sch
.SUBCKT foldedcascode_nmos_withdummies AVSS IBIAS AVDD PLUS MINUS VOUT D_ENA
*.PININFO AVSS:I IBIAS:I AVDD:I PLUS:I MINUS:I VOUT:O D_ENA:I
M23 IBIAS net3 AVSS AVSS sg13_lv_nmos w=8.5u l=5u ng=4 m=1
M25 IBIAS net2 net3 AVSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
M24 net10 net3 AVSS AVSS sg13_lv_nmos w=8.5u l=5u ng=4 m=1
M11 net10 net5 net4 AVDD sg13_lv_pmos w=14u l=2u ng=4 m=1
M12 net4 net4 AVDD AVDD sg13_lv_pmos w=14u l=2u ng=4 m=1
M18 AVSS net5 net8 AVDD sg13_lv_pmos w=14u l=0.5u ng=4 m=1
M17 net8 net4 AVDD AVDD sg13_lv_pmos w=14u l=2u ng=4 m=1
M9 net7 net4 AVDD AVDD sg13_lv_pmos w=14u l=2u ng=4 m=1
M5 net5 net8 net7 AVDD sg13_lv_pmos w=14u l=2u ng=4 m=1
M7 net5 net15 net6 AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
M3 net6 net5 AVSS AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
M30 net9 net3 AVSS AVSS sg13_lv_nmos w=8.5u l=5u ng=4 m=1
M1 net7 PLUS net9 AVSS sg13_lv_nmos w=6u l=1u ng=2 m=1
M2 net11 MINUS net9 AVSS sg13_lv_nmos w=6u l=1u ng=2 m=1
M42 AVDD net4 AVDD AVDD sg13_lv_pmos w=12u l=1u ng=4 m=1
M41 AVDD net8 AVDD AVDD sg13_lv_pmos w=12u l=1u ng=4 m=1
M38 AVSS net3 AVSS AVSS sg13_lv_nmos w=8u l=1u ng=4 m=1
M19 net1 D_ENA AVDD AVDD sg13_lv_pmos w=1u l=0.13u ng=1 m=1
M21 net2 net1 AVDD AVDD sg13_lv_pmos w=1u l=0.13u ng=1 m=1
M20 net1 D_ENA AVSS AVSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
M22 net2 net1 AVSS AVSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
M37 net11 AVSS AVSS AVSS sg13_lv_nmos w=6u l=1u ng=2 m=1
M6 VOUT net8 net11 AVDD sg13_lv_pmos w=14u l=2u ng=4 m=1
M0 net11 net4 AVDD AVDD sg13_lv_pmos w=14u l=2u ng=4 m=1
M8 VOUT net15 net12 AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
M4 net12 net5 AVSS AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
M29 net12 AVSS AVSS AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
M28 VOUT AVSS AVSS AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
M32 net11 AVDD AVDD AVDD sg13_lv_pmos w=14u l=2u ng=4 m=1
M33 VOUT AVDD AVDD AVDD sg13_lv_pmos w=7u l=2u ng=2 m=1
M13 net13 net4 AVDD AVDD sg13_lv_pmos w=14u l=2u ng=4 m=1
M15 net13 VOUT net14 AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
M16 net14 net14 AVSS AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
M14 net15 net14 AVSS AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
M10 AVDD VOUT net15 AVSS sg13_lv_nmos w=15u l=0.5u ng=4 m=1
M40 AVSS net15 AVSS AVSS sg13_lv_nmos w=8u l=1u ng=4 m=1
M39 net5 net1 AVSS AVSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
M36 net7 AVSS AVSS AVSS sg13_lv_nmos w=6u l=1u ng=2 m=1
M34 net5 AVDD AVDD AVDD sg13_lv_pmos w=7u l=2u ng=2 m=1
M27 net6 AVSS AVSS AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
M26 net5 AVSS AVSS AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
M35 net4 AVDD AVDD AVDD sg13_lv_pmos w=7u l=2u ng=2 m=1
M31 net14 AVSS AVSS AVSS sg13_lv_nmos w=3u l=2u ng=2 m=1
.ENDS
