<<<<<<< HEAD
** sch_path: /foss/designs/Thesis/workspace/thesis_hp/Schematics/Analog_Inverter/testbenches_Analog_Inverter/tb_Analog_Inverter_dc.sch
**.subckt tb_Analog_Inverter_dc
Vdd1 Vdd GND 1.5
Vss1 Vss GND 0
x1 Vdd v_in v_out Vss Analog_Inverter
Vin v_in GND dc 0 pulse(0 1.5 0 1n 1n 4n 10n)
=======
** sch_path: /foss/designs/thesis/workspace/thesis_hp/Designs/Analog_Inverter/Schematics/testbenches_Analog_Inverter/tb_Analog_Inverter_dc.sch
**.subckt tb_Analog_Inverter_dc
Vdd1 Vdd GND 1.5
Vss1 Vss GND 0
Vin v_in GND dc 0 pulse(0 1.5 0 1n 1n 4n 10n)
C1 v_out GND 50f m=1
x1 Vdd v_in v_out Vss Analog_Inverter
>>>>>>> f16623861683ae9920a8a8a8aa8d5da90f8a8425
**** begin user architecture code


*Vin v_in 0 dc 0 pulse(0 1.5 0 1n 1n 4n 10n)

.control
reset
dc vin 0 1.5 0.01
save all
let VP = 1.5
let vo_mid = VP/2
let dvout = deriv(v(v_out))
meas DC VSW find v(v_in) when v(v_out)=vo_mid
meas DC VIL find v(v_in) WHEN dvout=-1 CROSS=1
meas DC VIH find v(v_in) WHEN dvout=-1 CROSS=2
meas DC VOL find v(v_out) WHEN dvout=-1 CROSS=2
meas DC VOH find v(v_out) WHEN dvout=-1 CROSS=1
echo VTC measurements
print VSW
print VIL
print VIH
print VOH
print VOL
echo
*set filetype=binary
<<<<<<< HEAD
*write ./Analog_Inverter/simulations/tb_inv_dc.raw

plot v(v_out)
=======
write /designs/thesis/workspace/thesis_hp/designs/analog_inverter/schematics/simulations/tb_inv_dc.raw

plot v(v_out)
plot v(dvout)
>>>>>>> f16623861683ae9920a8a8a8aa8d5da90f8a8425


.endc
.end


 .lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends

<<<<<<< HEAD
* expanding   symbol:  /foss/designs/Thesis/workspace/thesis_hp/Schematics/Analog_Inverter/Analog_Inverter.sym # of pins=4
** sym_path: /foss/designs/Thesis/workspace/thesis_hp/Schematics/Analog_Inverter/Analog_Inverter.sym
** sch_path: /foss/designs/Thesis/workspace/thesis_hp/Schematics/Analog_Inverter/Analog_Inverter.sch
=======
* expanding   symbol:  /foss/designs/Thesis/workspace/thesis_hp/Designs/Analog_Inverter/Schematics/Analog_Inverter.sym # of pins=4
** sym_path: /foss/designs/Thesis/workspace/thesis_hp/Designs/Analog_Inverter/Schematics/Analog_Inverter.sym
** sch_path: /foss/designs/Thesis/workspace/thesis_hp/Designs/Analog_Inverter/Schematics/Analog_Inverter.sch
>>>>>>> f16623861683ae9920a8a8a8aa8d5da90f8a8425
.subckt Analog_Inverter vdd vin vout vss
*.ipin vin
*.iopin vdd
*.iopin vss
*.opin vout
<<<<<<< HEAD
XM1 vout vin vdd vdd sg13_lv_pmos w=40u l=0.52u ng=1 m=1
XM2 vout vin vss vss sg13_lv_nmos w=20u l=0.52u ng=1 m=1
=======
XM1 vout vin vdd vdd sg13_lv_pmos w=2u l=0.15u ng=1 m=1
XM2 vout vin vss vss sg13_lv_nmos w=1u l=0.15u ng=1 m=1
>>>>>>> f16623861683ae9920a8a8a8aa8d5da90f8a8425
.ends

.GLOBAL GND
.end
