.subckt FMD_QNC_ota_final_decoup VDD VSS
.ends
.end
