** sch_path: /foss/designs/thesis/workspace/thesis_hp/designs/otas/foldedcascode_nmos.sch
.subckt foldedcascode_nmos AVDD PLUS MINUS Vout Ibias AVSS
*.PININFO PLUS:I MINUS:I Vout:O AVDD:I AVSS:I Ibias:I
XM6 net5 PLUS net1 AVSS sg13_lv_nmos w=5u l=1u ng=1 m=1
XM8 net1 Ibias AVSS AVSS sg13_lv_nmos w=25u l=5u ng=3 m=1
XM21 net3 net4 AVSS AVSS sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM22 net2 net4 AVSS AVSS sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM7 net6 MINUS net1 AVSS sg13_lv_nmos w=5u l=1u ng=1 m=1
XM23 net4 net9 net2 AVSS sg13_lv_nmos w=1.5u l=0.5u ng=1 m=1
XM24 Vout net9 net3 AVSS sg13_lv_nmos w=1.5u l=0.5u ng=1 m=1
XM25 net4 net8 net5 AVDD sg13_lv_pmos w=6u l=0.5u ng=1 m=1
XM26 net5 net7 AVDD AVDD sg13_lv_pmos w=6u l=0.5u ng=1 m=1
XM27 Vout net8 net6 AVDD sg13_lv_pmos w=6u l=0.5u ng=1 m=1
XM28 net6 net7 AVDD AVDD sg13_lv_pmos w=6u l=0.5u ng=1 m=1
XM1 Ibias Ibias AVSS AVSS sg13_lv_nmos w=18u l=5u ng=2 m=1
XM2 net8 net8 net7 AVDD sg13_lv_pmos w=6u l=0.5u ng=2 m=1
XM3 net7 net7 AVDD AVDD sg13_lv_pmos w=6u l=0.5u ng=2 m=1
XM4 net9 net7 AVDD AVDD sg13_lv_pmos w=6u l=0.5u ng=2 m=1
XM5 net9 net9 AVSS AVSS sg13_lv_nmos w=1.5u l=0.5u ng=1 m=1
XM9 net8 Ibias AVSS AVSS sg13_lv_nmos w=25u l=5u ng=3 m=1
.ends
