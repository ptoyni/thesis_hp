* NGSPICE file created from FMD_QNC_ota_final_decoup.ext - technology: ihp-sg13g2

.subckt FMD_QNC_ota_decoup AVDD IBIAS VOUT MINUS PLUS AVSS
X0 a_n71700_n71833# a_n71700_n71833# a_n2191_3729# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X1 a_n2997_1502# a_n2191_3729# a_n7496_n2395# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X2 a_n71700_n71833# a_n36679_n4028# a_n7496_n1298# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X3 a_492_n6342# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X4 dw_n3357_1102# a_n2997_1502# a_n2227_3805# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X5 a_n2997_1502# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X6 a_n7496_n2395# a_n2191_3729# a_n2997_1502# dw_n3357_1102# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X7 a_n71700_n71833# a_n71700_n71833# a_n686_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X8 a_n2227_3805# a_n2191_3729# a_n71700_n71833# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=0.5u
X9 dw_n3357_1102# a_n2227_3805# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=1.02p pd=6.68u as=6.33942n ps=2.35229m w=3u l=0.5u
X10 a_n7496_n1298# a_n238_240# a_n2191_4205# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X11 a_10178_n5569# a_492_n4328# a_10269_2986# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X12 a_n71700_n71833# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.38p pd=2.38u as=9.72627n ps=3.82212m w=2u l=1u
X13 a_n722_n4252# a_10178_n5569# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X14 a_n2227_3805# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X15 dw_n3357_1102# a_n2997_1502# a_n2343_7081# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X16 dw_n3357_1102# a_n2997_1502# a_n2343_7081# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X17 a_n71700_n71833# a_n722_n4252# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.38p pd=2.38u as=0 ps=0 w=2u l=1u
X18 a_n2343_7081# a_n238_n912# a_n7496_n1298# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X19 dw_n3357_1102# a_n2227_3805# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=0.5u
X20 a_492_n4328# a_n71700_n71833# cap_cmim l=25.82u w=25.82u
X21 a_n686_n6342# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X22 a_n71700_n71833# a_n722_n4252# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.68p pd=4.68u as=0 ps=0 w=2u l=1u
X23 dw_n3357_1102# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=0.5u
X24 a_n2227_3805# a_n2191_3729# a_n71700_n71833# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=0.5u
X25 a_n7496_n1298# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X26 dw_n3357_1102# a_492_n4328# a_n722_n4252# a_n71700_n71833# sg13_lv_nmos ad=0.7125p pd=4.13u as=0.7125p ps=4.13u w=3.75u l=0.5u
X27 dw_n3357_1102# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=0.5u
X28 a_n2343_7081# a_n2227_3805# a_492_n4328# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X29 a_n7496_n1298# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X30 a_n2191_4205# a_n2227_3805# a_n2191_3729# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X31 a_n2191_3729# a_n2227_3805# a_n2191_4205# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X32 a_n71700_n71833# a_n36679_n4028# a_n7496_n2395# a_n71700_n71833# sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X33 a_n2343_7081# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X34 dw_n3357_1102# dw_n3357_1102# a_n2343_7081# dw_n3357_1102# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X35 a_n2343_7081# dw_n3357_1102# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X36 a_n71700_n71833# a_n36679_n4028# a_n36679_n4028# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X37 a_n71700_n71833# a_n2191_3729# a_492_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X38 dw_n3357_1102# a_n2997_1502# a_10269_2986# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X39 a_492_n6342# a_n722_n4252# a_492_n4328# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X40 dw_n3357_1102# a_n2997_1502# a_n2191_4205# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X41 a_n71700_n71833# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.38p pd=2.38u as=0 ps=0 w=2u l=1u
X42 a_10178_n5569# a_10178_n5569# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X43 dw_n3357_1102# a_n2227_3805# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=0.5u
X44 a_492_n4328# dw_n3357_1102# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X45 a_n2191_4205# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X46 a_n2343_7081# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=1.02p ps=6.68u w=3u l=1u
X47 dw_n3357_1102# a_n2997_1502# a_n2997_1502# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X48 a_n2191_3729# a_n2227_3805# a_n2191_4205# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X49 a_10269_2986# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X50 a_n71700_n71833# a_n2191_3729# a_n686_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X51 a_n36679_n4028# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X52 a_n2997_1502# a_n2191_3729# a_n7496_n2395# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X53 a_n71700_n71833# a_10178_n5569# a_n722_n4252# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X54 a_n686_n6342# a_n722_n4252# a_n2191_3729# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X55 dw_n3357_1102# a_n2997_1502# a_n2997_1502# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X56 a_n2191_4205# a_n238_240# a_n7496_n1298# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X57 a_n7496_n1298# a_n238_n912# a_n2343_7081# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X58 a_n36679_n4028# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X59 a_n722_n4252# a_492_n4328# dw_n3357_1102# a_n71700_n71833# sg13_lv_nmos ad=0.7125p pd=4.13u as=1.275p ps=8.18u w=3.75u l=0.5u
X60 a_492_n6342# a_n2191_3729# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X61 a_10269_2986# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X62 a_n2191_3729# dw_n3357_1102# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X63 a_10269_2986# a_492_n4328# a_10178_n5569# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X64 a_n722_n4252# a_492_n4328# dw_n3357_1102# a_n71700_n71833# sg13_lv_nmos ad=0.7125p pd=4.13u as=0.7125p ps=4.13u w=3.75u l=0.5u
X65 a_492_n4328# a_n722_n4252# a_492_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X66 a_10178_n5569# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X67 a_n2997_1502# dw_n3357_1102# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X68 a_n2227_3805# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X69 a_n2343_7081# dw_n3357_1102# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X70 a_n71700_n71833# a_n36679_n4028# a_n7496_n1298# a_n71700_n71833# sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X71 a_n71700_n71833# a_n36679_n4028# a_n7496_n2395# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X72 a_n2191_4205# a_n2227_3805# a_n2191_3729# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X73 a_n71700_n71833# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.38p pd=2.38u as=0 ps=0 w=2u l=1u
X74 a_n71700_n71833# a_n71700_n71833# a_n2343_7081# a_n71700_n71833# sg13_lv_nmos ad=1.02p pd=6.68u as=0.57p ps=3.38u w=3u l=1u
X75 a_n71700_n71833# a_n2191_3729# a_n2227_3805# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=0.5u
X76 dw_n3357_1102# dw_n3357_1102# a_492_n4328# dw_n3357_1102# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X77 a_n686_n6342# a_n2191_3729# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X78 a_n2191_3729# a_n722_n4252# a_n686_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X79 a_n2343_7081# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X80 dw_n3357_1102# a_n2227_3805# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=0.5u
X81 a_n2997_1502# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X82 a_n71700_n71833# a_n71700_n71833# a_10178_n5569# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X83 a_n71700_n71833# a_n722_n4252# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.38p pd=2.38u as=0 ps=0 w=2u l=1u
X84 a_n71700_n71833# a_n71700_n71833# a_n2191_4205# a_n71700_n71833# sg13_lv_nmos ad=1.02p pd=6.68u as=0.57p ps=3.38u w=3u l=1u
X85 dw_n3357_1102# a_n2997_1502# a_n2191_4205# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X86 a_492_n4328# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X87 a_n71700_n71833# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.68p pd=4.68u as=0 ps=0 w=2u l=1u
X88 dw_n3357_1102# dw_n3357_1102# a_n2997_1502# dw_n3357_1102# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X89 a_n7496_n2395# a_n2191_3729# a_n2997_1502# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X90 a_n71700_n71833# a_n722_n4252# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.38p pd=2.38u as=0 ps=0 w=2u l=1u
X91 a_n2343_7081# a_n2227_3805# a_492_n4328# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X92 a_492_n4328# a_n2227_3805# a_n2343_7081# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X93 a_n7496_n2395# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X94 dw_n3357_1102# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.57p pd=3.38u as=0 ps=0 w=3u l=0.5u
X95 dw_n3357_1102# dw_n3357_1102# a_n2191_3729# dw_n3357_1102# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X96 a_n71700_n71833# a_n71700_n71833# a_492_n4328# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X97 dw_n3357_1102# a_n2997_1502# a_10269_2986# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X98 dw_n3357_1102# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=1.02p pd=6.68u as=0 ps=0 w=3u l=0.5u
X99 a_n7496_n2395# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X100 dw_n3357_1102# dw_n3357_1102# a_n2343_7081# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X101 a_n71700_n71833# a_10178_n5569# a_10178_n5569# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X102 a_n71700_n71833# a_n71700_n71833# a_492_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X103 dw_n3357_1102# a_n2997_1502# a_n2227_3805# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X104 a_n2191_3729# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X105 a_n71700_n71833# a_n36679_n4028# a_n36679_n4028# a_n71700_n71833# sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X106 a_n2191_4205# a_n2997_1502# dw_n3357_1102# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X107 a_n71700_n71833# a_n2191_3729# a_n2227_3805# dw_n3357_1102# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=0.5u
X108 a_n2191_4205# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=1.02p ps=6.68u w=3u l=1u
X109 dw_n3357_1102# a_492_n4328# a_n722_n4252# a_n71700_n71833# sg13_lv_nmos ad=1.275p pd=8.18u as=0.7125p ps=4.13u w=3.75u l=0.5u
X110 a_492_n4328# a_n2227_3805# a_n2343_7081# dw_n3357_1102# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
.ends
