.subckt foldedcascode_nmos_withdummies VDD VSS
.ends
.end
