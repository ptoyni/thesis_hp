.subckt complete_schematic_pads VDD VSS
.ends
.end
