* Extracted by KLayout with SG13G2 LVS runset on : 12/07/2025 23:28

.SUBCKT ota_final AVSS PLUS AVDD VOUT IBIAS MINUS
M$1 AVDD VOUT \$18333 AVSS sg13_lv_nmos L=0.5u W=15u AS=3.4125p AD=3.4125p
+ PS=20.57u PD=20.57u
M$5 AVSS IBIAS IBIAS AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$9 AVSS IBIAS \$19330 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$13 AVSS IBIAS \$19329 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$17 AVSS AVSS \$19441 AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$18 \$19441 MINUS \$19329 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p
+ PS=6.76u PD=6.76u
M$19 \$19329 PLUS \$19657 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p
+ PS=6.76u PD=6.76u
M$20 \$19657 AVSS AVSS AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$25 \$19330 \$18830 \$19331 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
M$29 AVSS \$18830 \$19333 AVDD sg13_lv_pmos L=0.5u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
M$33 \$18334 VOUT \$18335 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$35 AVSS AVSS \$18334 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$36 \$18334 \$18334 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$37 AVSS \$18334 \$18333 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$41 AVSS AVSS VOUT AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$42 VOUT \$18333 \$I481451 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$45 AVSS AVSS \$I481450 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$46 \$I481450 \$18830 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$49 AVSS AVSS \$I481451 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$50 \$I481451 \$18830 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$53 AVSS AVSS \$18830 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$54 \$18830 \$18333 \$I481450 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$57 AVDD AVDD \$19331 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p
+ PS=11.56u PD=11.56u
M$58 \$19331 \$19331 AVDD AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$59 AVDD \$19331 \$19333 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$61 AVDD \$19331 \$18335 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$71 AVDD AVDD \$18830 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p
+ PS=11.56u PD=11.56u
M$72 \$18830 \$19333 \$19657 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$77 AVDD AVDD VOUT AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$78 VOUT \$19333 \$19441 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$83 AVDD AVDD \$19441 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
M$85 AVDD \$19331 \$19657 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$87 AVDD \$19331 \$19441 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
.ENDS ota_final
