* NGSPICE file created from FMD_QNC_ota_final_esd.ext - technology: ihp-sg13g2

.subckt FMD_QNC_ota_final_esd IBIAS MINUS PLUS VOUT AVDD AVSS
X0 a_n1791_7045# a_n1791_7045# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X1 dw_n3357_2616# a_n1791_7045# a_n2227_3805# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X2 a_n71700_n71833# a_n36679_n4028# a_n7496_n1298# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X3 a_n1791_7045# a_n2191_3729# a_n7496_n2395# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X4 a_n71700_n71833# a_n71700_n71833# a_n2191_3729# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X5 a_492_n6342# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X6 a_n7496_n2395# a_n2191_3729# a_n1791_7045# dw_n3357_2616# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X7 a_n2227_3805# a_n2191_3729# a_n71700_n71833# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=0.5u
X8 a_n71700_n71833# a_n71700_n71833# a_n686_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X9 a_n7496_n1298# a_n238_240# a_n2191_4205# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X10 a_10178_n5569# a_492_n4328# a_10269_2986# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X11 a_n2227_3805# a_n1791_7045# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X12 a_n722_n4252# a_10178_n5569# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X13 dw_n3357_2616# a_n1791_7045# a_n2343_7081# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X14 dw_n3357_2616# a_n1791_7045# a_n2343_7081# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X15 a_n2343_7081# a_n238_n912# a_n7496_n1298# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X16 a_n686_n6342# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X17 a_492_n4328# a_n71700_n71833# cap_cmim l=25.82u w=25.82u
X18 a_n7496_n1298# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X19 a_n2227_3805# a_n2191_3729# a_n71700_n71833# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=0.5u
X20 dw_n3357_2616# a_492_n4328# a_n722_n4252# a_n71700_n71833# sg13_lv_nmos ad=0.7125p pd=4.13u as=0.7125p ps=4.13u w=3.75u l=0.5u
X21 a_n2343_7081# a_n2227_3805# a_492_n4328# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X22 a_n7496_n1298# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X23 a_n2343_7081# a_n1791_7045# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X24 dw_n3357_2616# dw_n3357_2616# a_n2343_7081# dw_n3357_2616# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X25 a_n2191_3729# a_n2227_3805# a_n2191_4205# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X26 a_n2191_4205# a_n2227_3805# a_n2191_3729# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X27 a_n71700_n71833# a_n36679_n4028# a_n7496_n2395# a_n71700_n71833# sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X28 a_n2343_7081# dw_n3357_2616# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X29 dw_n3357_2616# a_n1791_7045# a_10269_2986# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X30 a_n71700_n71833# a_n36679_n4028# a_n36679_n4028# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X31 a_n71700_n71833# a_n2191_3729# a_492_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X32 a_492_n6342# a_n722_n4252# a_492_n4328# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X33 dw_n3357_2616# a_n1791_7045# a_n2191_4205# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X34 a_10178_n5569# a_10178_n5569# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X35 a_n2191_4205# a_n1791_7045# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X36 a_492_n4328# dw_n3357_2616# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X37 a_n2191_3729# a_n2227_3805# a_n2191_4205# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X38 a_10269_2986# a_n1791_7045# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X39 dw_n3357_2616# a_n1791_7045# a_n1791_7045# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X40 a_n2343_7081# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=1.02p ps=6.68u w=3u l=1u
X41 a_n71700_n71833# a_n2191_3729# a_n686_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X42 dw_n3357_2616# a_n1791_7045# a_n1791_7045# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X43 a_n1791_7045# a_n2191_3729# a_n7496_n2395# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X44 a_n36679_n4028# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X45 a_n686_n6342# a_n722_n4252# a_n2191_3729# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X46 a_n71700_n71833# a_10178_n5569# a_n722_n4252# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X47 a_n7496_n1298# a_n238_n912# a_n2343_7081# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X48 a_n2191_4205# a_n238_240# a_n7496_n1298# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X49 a_n36679_n4028# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X50 a_n2191_3729# dw_n3357_2616# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X51 a_10269_2986# a_n1791_7045# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X52 a_492_n4328# a_n722_n4252# a_492_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X53 a_492_n6342# a_n2191_3729# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X54 a_n722_n4252# a_492_n4328# dw_n3357_2616# a_n71700_n71833# sg13_lv_nmos ad=0.7125p pd=4.13u as=0.7125p ps=4.13u w=3.75u l=0.5u
X55 a_n722_n4252# a_492_n4328# dw_n3357_2616# a_n71700_n71833# sg13_lv_nmos ad=0.7125p pd=4.13u as=1.275p ps=8.18u w=3.75u l=0.5u
X56 a_10269_2986# a_492_n4328# a_10178_n5569# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X57 a_10178_n5569# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X58 a_n2343_7081# dw_n3357_2616# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X59 a_n2227_3805# a_n1791_7045# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X60 a_n1791_7045# dw_n3357_2616# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X61 a_n71700_n71833# a_n36679_n4028# a_n7496_n1298# a_n71700_n71833# sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X62 a_n71700_n71833# a_n36679_n4028# a_n7496_n2395# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X63 a_n2191_4205# a_n2227_3805# a_n2191_3729# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X64 a_n71700_n71833# a_n71700_n71833# a_n2343_7081# a_n71700_n71833# sg13_lv_nmos ad=1.02p pd=6.68u as=0.57p ps=3.38u w=3u l=1u
X65 dw_n3357_2616# dw_n3357_2616# a_492_n4328# dw_n3357_2616# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X66 a_n71700_n71833# a_n2191_3729# a_n2227_3805# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=0.5u
X67 a_n2191_3729# a_n722_n4252# a_n686_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X68 a_n686_n6342# a_n2191_3729# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X69 dw_n3357_2616# a_n1791_7045# a_n2191_4205# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X70 a_n2343_7081# a_n1791_7045# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X71 dw_n3357_2616# dw_n3357_2616# a_n1791_7045# dw_n3357_2616# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X72 a_n1791_7045# a_n1791_7045# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X73 a_n71700_n71833# a_n71700_n71833# a_n2191_4205# a_n71700_n71833# sg13_lv_nmos ad=1.02p pd=6.68u as=0.57p ps=3.38u w=3u l=1u
X74 a_492_n4328# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X75 a_n71700_n71833# a_n71700_n71833# a_10178_n5569# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X76 a_492_n4328# a_n2227_3805# a_n2343_7081# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X77 a_n2343_7081# a_n2227_3805# a_492_n4328# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X78 a_n7496_n2395# a_n2191_3729# a_n1791_7045# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X79 a_n7496_n2395# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X80 dw_n3357_2616# dw_n3357_2616# a_n2191_3729# dw_n3357_2616# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X81 dw_n3357_2616# a_n1791_7045# a_10269_2986# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X82 a_n71700_n71833# a_n71700_n71833# a_492_n4328# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X83 dw_n3357_2616# dw_n3357_2616# a_n2343_7081# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X84 dw_n3357_2616# a_n1791_7045# a_n2227_3805# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X85 a_n7496_n2395# a_n36679_n4028# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X86 a_n71700_n71833# a_n36679_n4028# a_n36679_n4028# a_n71700_n71833# sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X87 a_n2191_3729# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X88 a_n71700_n71833# a_n71700_n71833# a_492_n6342# a_n71700_n71833# sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X89 a_n71700_n71833# a_10178_n5569# a_10178_n5569# a_n71700_n71833# sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X90 a_n2191_4205# a_n1791_7045# dw_n3357_2616# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X91 a_n71700_n71833# a_n2191_3729# a_n2227_3805# dw_n3357_2616# sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=0.5u
X92 a_492_n4328# a_n2227_3805# a_n2343_7081# dw_n3357_2616# sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X93 a_n2191_4205# a_n71700_n71833# a_n71700_n71833# a_n71700_n71833# sg13_lv_nmos ad=0.57p pd=3.38u as=1.02p ps=6.68u w=3u l=1u
X94 dw_n3357_2616# a_492_n4328# a_n722_n4252# a_n71700_n71833# sg13_lv_nmos ad=1.275p pd=8.18u as=0.7125p ps=4.13u w=3.75u l=0.5u
C0 a_n7496_n2395# a_n2227_3805# 0.05824f
C1 a_n1791_7045# a_n2343_7081# 1.2779f
C2 a_n238_n912# a_n7496_n1298# 0.26247f
C3 a_n238_n912# a_n2191_3729# 0.10776f
C4 a_n7496_n2395# a_492_n4328# 0.2268f
C5 dw_n3357_2616# w_9484_45# 0.03598f
C6 a_n238_n912# a_n2191_4205# 0.14151f
C7 dw_n3357_2616# a_n238_240# 2.00834f
C8 m3_n71700_n71833# m4_n71700_n71833# 0.39453p
C9 a_10269_2986# a_n2227_3805# 0.1057f
C10 a_n2343_7081# a_n7496_n2395# 0.0628f
C11 dw_n3357_2616# m1_n6131_n62493# 0.22767f
C12 a_492_n4328# a_10269_2986# 0.69235f
C13 m7_n71700_n71833# m6_n71120_n71253# 49.114f
C14 a_n1791_7045# a_n7496_n2395# 0.25761f
C15 m6_n71700_n71833# m7_n71700_n71833# 76.089f
C16 a_n2191_3729# a_n2227_3805# 1.43394f
C17 a_n2191_3729# a_n686_n6342# 0.43014f
C18 dw_n3357_2616# a_n238_n912# 2.08158f
C19 m6_n71700_n71833# m5_n71700_n71833# 0.25064p
C20 a_492_n4328# a_n2191_3729# 0.28555f
C21 a_n63343_11041# m1_n64157_14354# 0.24502p
C22 a_n1791_7045# a_10269_2986# 0.8497f
C23 a_n2227_3805# a_n2191_4205# 1.02301f
C24 a_n238_240# a_n238_n912# 0.09545f
C25 a_n722_n4252# a_n2191_3729# 0.3829f
C26 a_n2343_7081# a_n7496_n1298# 0.25316f
C27 a_n7496_n2395# a_n36679_n4028# 1.35216f
C28 m2_n71700_n71833# m3_n71700_n71833# 0.39453p
C29 a_n1791_7045# a_n2191_3729# 0.95025f
C30 a_n5317_n65806# m1_n6131_n62493# 0.24502p
C31 a_n2343_7081# a_n2191_4205# 0.42257f
C32 dw_n3357_2616# w_9059_n1941# 0.02677f
C33 m1_n6133_51337# a_n5319_48024# 0.24502p
C34 m3_n71262_n71395# m2_n71262_n71395# 0.39413p
C35 a_n1791_7045# a_n2191_4205# 0.95151f
C36 dw_n3357_2616# a_n2227_3805# 11.6462f
C37 a_52706_n30940# m1_51892_n27627# 0.24502p
C38 a_n7496_n2395# a_n7496_n1298# 0.0392f
C39 dw_n3357_2616# a_492_n4328# 5.09315f
C40 a_n7496_n2395# a_n2191_3729# 1.18183f
C41 a_n238_240# a_n2227_3805# 0.58224f
C42 dw_n3357_2616# w_n3357_2616# 0.04671f
C43 a_492_n4328# a_10178_n5569# 0.33532f
C44 a_n238_240# a_492_n4328# 0.06043f
C45 a_n7496_n2395# a_n2191_4205# 0.0626f
C46 dw_n3357_2616# a_n722_n4252# 0.94287f
C47 dw_n3357_2616# a_n2343_7081# 3.59868f
C48 a_n7496_n1298# a_n36679_n4028# 1.39083f
C49 a_n2191_3729# a_n36679_n4028# 0.39006f
C50 a_n2191_3729# a_10269_2986# 0.01919f
C51 a_492_n4328# a_492_n6342# 0.11125f
C52 a_n1791_7045# dw_n3357_2616# 26.2822f
C53 a_n47332_n65813# m1_n48146_n62500# 0.24502p
C54 m3_n71262_n71395# m4_n71262_n71395# 0.39413p
C55 a_n722_n4252# a_10178_n5569# 0.27513f
C56 a_n238_240# a_n2343_7081# 0.12558f
C57 a_n1791_7045# a_n238_240# 0.55923f
C58 m5_n71216_n71349# m6_n71120_n71253# 0.16179p
C59 a_n722_n4252# a_492_n6342# 0.26872f
C60 a_n2191_3729# a_n7496_n1298# 0.10311f
C61 dw_n3357_2616# a_n7496_n2395# 2.16832f
C62 dw_n3357_2616# a_15657_n65815# 0.24502p
C63 a_n7496_n1298# a_n2191_4205# 0.31895f
C64 a_n2191_3729# a_n2191_4205# 0.26032f
C65 a_n238_240# a_n7496_n2395# 0.57854f
C66 a_n2343_7081# a_n238_n912# 0.26338f
C67 dw_n3357_2616# a_n36679_n4028# 16.5402f
C68 a_n63359_n30959# m1_n64173_n27646# 0.24502p
C69 dw_n3357_2616# a_10269_2986# 1.32667f
C70 a_36679_48076# m1_35865_51389# 0.24502p
C71 m2_n71700_n71833# m1_n71700_n71833# 0.39453p
C72 a_36681_n65774# m1_35867_n62461# 0.24502p
C73 a_10269_2986# a_10178_n5569# 0.11798f
C74 a_492_n4328# a_n2227_3805# 0.99098f
C75 a_52655_11010# m1_51841_14323# 0.24502p
C76 dw_n3357_2616# a_n2191_3729# 7.13697f
C77 a_n7496_n2395# a_n238_n912# 0.05813f
C78 a_n238_240# a_n7496_n1298# 0.36761f
C79 a_n238_240# a_n2191_3729# 0.12975f
C80 a_n2343_7081# a_n2227_3805# 1.09777f
C81 m1_n71262_n71395# m2_n71262_n71395# 0.39413p
C82 a_n722_n4252# a_n686_n6342# 0.24377f
C83 dw_n3357_2616# a_n2191_4205# 2.18016f
C84 a_n722_n4252# a_492_n4328# 1.47142f
C85 m1_n48145_51360# a_n47331_48047# 0.24502p
C86 a_n238_n912# a_n36679_n4028# 0.13883f
C87 a_n2343_7081# a_492_n4328# 0.25886f
C88 a_n1791_7045# a_n2227_3805# 1.27969f
C89 a_n2191_3729# a_492_n6342# 0.2849f
C90 m5_n71700_n71833# m4_n71700_n71833# 0.39453p
C91 m4_n71262_n71395# m5_n71216_n71349# 0.34892p
C92 a_n238_240# a_n2191_4205# 0.29063f
C93 m7_14896_51462# a_n71700_n71833# 17.8454f $ **FLOATING
C94 m7_n27115_51490# a_n71700_n71833# 17.8453f $ **FLOATING
C95 m7_n71700_n71833# a_n71700_n71833# 0.19092p
C96 m6_n71120_n71253# a_n71700_n71833# 0.21787p
C97 m6_n71700_n71833# a_n71700_n71833# 0.21939p
C98 m5_n71216_n71349# a_n71700_n71833# 0.16053p
C99 m5_n71700_n71833# a_n71700_n71833# 0.16155p
C100 m4_n71262_n71395# a_n71700_n71833# 0.16966p
C101 m4_n71700_n71833# a_n71700_n71833# 0.17068p
C102 m3_n71262_n71395# a_n71700_n71833# 0.1829p
C103 m3_n71700_n71833# a_n71700_n71833# 0.184p
C104 m2_n71262_n71395# a_n71700_n71833# 0.203p
C105 m2_n71700_n71833# a_n71700_n71833# 0.20422p
C106 m1_35867_n62461# a_n71700_n71833# 97.463f
C107 m1_n6131_n62493# a_n71700_n71833# 97.32021f
C108 m1_n48146_n62500# a_n71700_n71833# 97.63829f
C109 m1_51892_n27627# a_n71700_n71833# 98.1675f
C110 m1_n64173_n27646# a_n71700_n71833# 98.3161f
C111 m1_51895_n6638# a_n71700_n71833# 0.25703p $ **FLOATING
C112 m1_n64159_n6608# a_n71700_n71833# 0.25702p $ **FLOATING
C113 m1_51841_14323# a_n71700_n71833# 98.38451f
C114 m1_n64157_14354# a_n71700_n71833# 98.3119f
C115 m1_35865_51389# a_n71700_n71833# 99.30901f
C116 m1_n6133_51337# a_n71700_n71833# 84.1929f
C117 m1_n48145_51360# a_n71700_n71833# 99.4816f
C118 m1_n71262_n71395# a_n71700_n71833# 0.43621p
C119 m1_n71700_n71833# a_n71700_n71833# 0.43781p
C120 a_n26374_n65784# a_n71700_n71833# 0.24502p $ **FLOATING
C121 a_10178_n5569# a_n71700_n71833# 4.78595f $ **FLOATING
C122 a_492_n6342# a_n71700_n71833# 1.43265f $ **FLOATING
C123 a_n686_n6342# a_n71700_n71833# 1.39642f $ **FLOATING
C124 a_n722_n4252# a_n71700_n71833# 7.22686f $ **FLOATING
C125 a_n7496_n2395# a_n71700_n71833# 7.26254f $ **FLOATING
C126 a_n36679_n4028# a_n71700_n71833# 76.9817f $ **FLOATING
C127 a_n7496_n1298# a_n71700_n71833# 2.98906f $ **FLOATING
C128 a_n238_240# a_n71700_n71833# 56.1234f $ **FLOATING
C129 a_n238_n912# a_n71700_n71833# 54.7545f $ **FLOATING
C130 a_10269_2986# a_n71700_n71833# 4.11048f $ **FLOATING
C131 a_n2227_3805# a_n71700_n71833# 7.43891f $ **FLOATING
C132 a_492_n4328# a_n71700_n71833# 84.93761f $ **FLOATING
C133 a_n2191_3729# a_n71700_n71833# 16.4072f $ **FLOATING
C134 a_n2191_4205# a_n71700_n71833# 3.23251f $ **FLOATING
C135 a_n2343_7081# a_n71700_n71833# 2.53274f $ **FLOATING
C136 a_n1791_7045# a_n71700_n71833# 10.8306f $ **FLOATING
C137 dw_n3357_2616# a_n71700_n71833# 0.33596p $ **FLOATING
.ends
