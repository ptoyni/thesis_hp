* NGSPICE file created from ota_final.ext - technology: ihp-sg13g2

.subckt ota_final MINUS AVDD AVSS PLUS VOUT IBIAS
X0 AVSS IBIAS a_n7496_n1298# AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X1 AVSS AVSS a_n686_n3376# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X2 a_492_n6342# AVSS AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X3 a_7669_2986# a_n1791_7045# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X4 a_n1791_7045# a_n2191_3729# a_n7496_n2395# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X5 AVSS AVSS a_n686_n5390# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X6 a_n7496_n1298# PLUS a_n314_276# AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X7 a_7669_5842# a_n1791_7045# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X8 a_37_7081# a_n1791_7045# a_n439_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X9 a_1941_7081# a_n1791_7045# a_1465_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X10 a_n314_n876# MINUS a_n7496_n1298# AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X11 a_n722_n4252# VOUT AVDD AVSS sg13_lv_nmos ad=0.7125p pd=4.13u as=0.7125p ps=4.13u w=3.75u l=0.5u
X12 a_n722_n4252# VOUT AVDD AVSS sg13_lv_nmos ad=0.7125p pd=4.13u as=1.275p ps=8.18u w=3.75u l=0.5u
X13 a_7669_1082# AVDD AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X14 a_7578_n5569# AVSS AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X15 a_n686_n6342# AVSS AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X16 a_7669_3938# a_n1791_7045# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X17 a_n7496_n1298# IBIAS AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X18 AVSS a_n2191_3729# a_n2227_3805# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=0.5u
X19 AVDD AVDD a_7669_6794# AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X20 a_1623_5158# a_n2227_3805# a_1623_4682# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X21 a_n7496_n1298# IBIAS AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X22 AVSS AVSS a_7578_n5569# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X23 a_n439_7081# a_n1791_7045# a_n915_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X24 a_2893_7081# AVDD a_2417_7081# AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X25 a_n2191_4681# a_n2227_3805# a_n2191_4205# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X26 a_n2191_4205# a_n2227_3805# a_n2191_3729# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X27 AVSS IBIAS a_n7496_n2395# AVSS sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X28 a_n2343_7081# AVDD a_n2811_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X29 a_n7496_n2395# a_n2191_3729# a_n1791_7045# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X30 AVSS IBIAS IBIAS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X31 a_492_n5866# a_n2191_3729# a_492_n6342# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X32 AVDD a_n1791_7045# a_7669_4890# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X33 a_492_n3852# a_n722_n4252# a_492_n4328# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X34 AVDD a_n1791_7045# a_513_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X35 a_n1391_7081# a_n1791_7045# a_n1867_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X36 VOUT AVDD AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X37 AVDD a_n1791_7045# a_7669_2034# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X38 a_n1791_7045# a_n2191_3729# a_n7496_n2395# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X39 AVSS a_7578_n5569# a_7578_n5569# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X40 a_n2191_3729# a_n2227_3805# a_n2191_5157# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X41 a_n314_n876# AVSS AVSS AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=1.02p ps=6.68u w=3u l=1u
X42 a_n2227_3805# a_n2191_3729# AVSS AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=0.5u
X43 AVSS a_n2191_3729# a_n2227_3805# AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=0.5u
X44 a_n686_n5866# a_n2191_3729# a_n686_n6342# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X45 IBIAS IBIAS AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X46 a_n686_n3852# a_n722_n4252# a_n686_n4328# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X47 a_7578_n5569# VOUT a_9374_n4648# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X48 a_7669_6794# a_n1791_7045# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X49 AVDD a_n1791_7045# a_7669_5842# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X50 a_n7496_n1298# MINUS a_n314_n876# AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X51 a_n314_276# PLUS a_n7496_n1298# AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=0.57p ps=3.38u w=3u l=1u
X52 IBIAS IBIAS AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X53 a_8530_n5569# a_7578_n5569# AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X54 a_n2191_3729# AVDD AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=1.19p ps=7.68u w=3.5u l=2u
X55 a_n7496_n2395# a_n2191_3729# a_n1791_7045# AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X56 a_492_n3376# a_n722_n4252# a_492_n3852# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X57 a_492_n5390# a_n2191_3729# a_492_n5866# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X58 AVDD VOUT a_n722_n4252# AVSS sg13_lv_nmos ad=1.275p pd=8.18u as=0.7125p ps=4.13u w=3.75u l=0.5u
X59 a_2417_7081# AVDD a_1941_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X60 a_7669_2034# a_n1791_7045# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X61 AVSS IBIAS a_n7496_n1298# AVSS sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X62 AVSS IBIAS a_n7496_n2395# AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X63 a_n2191_5157# a_n2227_3805# a_n2191_4681# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X64 AVSS AVSS a_n314_n876# AVSS sg13_lv_nmos ad=1.02p pd=6.68u as=0.57p ps=3.38u w=3u l=1u
X65 AVDD AVDD VOUT AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X66 a_n2227_3805# a_n2191_3729# AVSS AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=0.5u
X67 a_n686_n3376# a_n722_n4252# a_n686_n3852# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X68 a_n686_n5390# a_n2191_3729# a_n686_n5866# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X69 a_n915_7081# a_n1791_7045# a_n1391_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X70 a_1465_7081# a_n1791_7045# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X71 AVSS AVSS a_n314_276# AVSS sg13_lv_nmos ad=1.02p pd=6.68u as=0.57p ps=3.38u w=3u l=1u
X72 a_492_n4328# AVSS AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X73 a_7578_n5569# a_7578_n5569# AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
X74 a_1623_4682# a_n2227_3805# a_1623_4206# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X75 a_1623_4206# a_n2227_3805# VOUT AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X76 AVDD a_n1791_7045# a_7669_2986# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X77 AVDD VOUT a_n722_n4252# AVSS sg13_lv_nmos ad=0.7125p pd=4.13u as=0.7125p ps=4.13u w=3.75u l=0.5u
X78 a_n7496_n2395# IBIAS AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.40375p ps=2.505u w=2.125u l=5u
X79 AVDD AVDD a_n2191_3729# AVDD sg13_lv_pmos ad=1.19p pd=7.68u as=0.665p ps=3.88u w=3.5u l=2u
X80 AVSS AVSS a_492_n3376# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X81 a_n1867_7081# AVDD a_n2343_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X82 AVDD a_n1791_7045# a_7669_1082# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X83 a_n7496_n2395# IBIAS AVSS AVSS sg13_lv_nmos ad=0.40375p pd=2.505u as=0.7225p ps=4.93u w=2.125u l=5u
X84 AVSS IBIAS IBIAS AVSS sg13_lv_nmos ad=0.7225p pd=4.93u as=0.40375p ps=2.505u w=2.125u l=5u
X85 a_n686_n4328# AVSS AVSS AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X86 AVSS AVSS a_492_n5390# AVSS sg13_lv_nmos ad=0.51p pd=3.68u as=0.285p ps=1.88u w=1.5u l=2u
X87 a_7669_4890# a_n1791_7045# AVDD AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X88 a_513_7081# a_n1791_7045# a_37_7081# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X89 a_9374_n4648# VOUT a_7578_n5569# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.51p ps=3.68u w=1.5u l=2u
X90 VOUT a_n2227_3805# a_1623_5158# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X91 AVDD a_n1791_7045# a_7669_3938# AVDD sg13_lv_pmos ad=0.665p pd=3.88u as=0.665p ps=3.88u w=3.5u l=2u
X92 a_n314_276# AVSS AVSS AVSS sg13_lv_nmos ad=0.57p pd=3.38u as=1.02p ps=6.68u w=3u l=1u
X93 AVSS a_7578_n5569# a_8530_n5569# AVSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.285p ps=1.88u w=1.5u l=2u
C0 a_n1391_7081# a_n314_276# 0.07138f
C1 a_51497_16180# VOUT 19.2483f
C2 a_n65951_36680# MINUS 19.7057f
C3 a_n314_276# a_n7496_n1298# 0.31866f
C4 a_n722_n4252# VOUT 1.05112f
C5 a_n2191_3729# m1_492_n6334# 0.28459f
C6 a_n2191_3729# PLUS 1.2526f
C7 a_n2227_3805# a_7669_2034# 0.07179f
C8 a_492_n4328# VOUT 0.03151f
C9 a_9374_n4648# VOUT 0.57151f
C10 a_n314_n876# VOUT 0.24724f
C11 a_n65932_15680# IBIAS 19.2326f
C12 a_n7496_n1298# a_n7496_n2395# 0.03162f
C13 a_n686_n3852# m1_n686_n6334# 0.03124f
C14 a_n722_n4252# m1_492_n6334# 0.30261f
C15 a_n314_276# a_n7496_n2395# 0.06208f
C16 a_n314_276# AVDD 1.50448f
C17 a_n686_n5390# m1_n686_n6334# 0.03177f
C18 a_n686_n6342# m1_n686_n6334# 0.03135f
C19 a_n314_n876# PLUS 0.11802f
C20 a_n7496_n2395# AVDD 1.59102f
C21 a_n7496_n1298# MINUS 0.26219f
C22 a_n65944_n47320# PLUS 19.9373f
C23 a_n314_276# MINUS 0.13825f
C24 a_1623_5158# a_n314_n876# 0.07222f
C25 m2_n77751_n74411# m3_n77751_n74411# 0.42115p
C26 m4_n77751_n74411# m5_n77705_n74365# 0.37285p
C27 a_n7496_n2395# MINUS 0.02524f
C28 a_n7496_n1298# IBIAS 1.39068f
C29 AVDD MINUS 2.03495f
C30 a_n65898_n5320# IBIAS 19.1558f
C31 a_7669_4890# a_9374_n4648# 0.06998f
C32 a_513_7081# a_n314_276# 0.07138f
C33 a_n439_7081# a_n314_n876# 0.07227f
C34 a_n2227_3805# a_n314_276# 1.01341f
C35 a_n2191_3729# a_n2191_4681# 0.07259f
C36 a_n2191_3729# a_n686_n3376# 0.03238f
C37 a_n2191_4205# a_n314_276# 0.07238f
C38 a_n7496_n2395# IBIAS 1.27464f
C39 m1_492_n6334# VOUT 0.10634f
C40 AVDD IBIAS 1.77558f
C41 a_n722_n4252# a_8530_n5569# 0.03137f
C42 m1_n77751_n74411# m2_n77751_n74411# 0.42115p
C43 a_n2227_3805# a_n7496_n2395# 0.04128f
C44 m2_n78189_n74849# m3_n78189_n74849# 0.42142p
C45 a_n2227_3805# AVDD 10.7658f
C46 m4_n78189_n74849# m5_n78189_n74849# 0.42142p
C47 a_37_7081# AVDD 0.07097f
C48 a_n1791_7045# a_n314_276# 0.9453f
C49 a_n2191_3729# a_n686_n4328# 0.03197f
C50 a_n2191_3729# a_n7496_n1298# 0.0862f
C51 MINUS IBIAS 0.13224f
C52 a_n2191_3729# a_n314_276# 0.24784f
C53 a_n1791_7045# a_7669_3938# 0.07097f
C54 a_n1791_7045# a_n7496_n2395# 0.25749f
C55 a_n1791_7045# AVDD 26.2642f
C56 a_n722_n4252# a_7578_n5569# 0.27873f
C57 a_n2191_3729# a_n7496_n2395# 1.17804f
C58 a_n2191_3729# AVDD 6.99442f
C59 w_n3276_2616# AVDD 0.08678f
C60 a_7578_n5569# a_9374_n4648# 0.11785f
C61 a_n7496_n1298# a_n314_n876# 0.25315f
C62 m1_n78189_n74849# m2_n78189_n74849# 0.42142p
C63 a_n49210_n62320# PLUS 19.9733f
C64 a_1623_4682# VOUT 0.07308f
C65 a_n314_276# a_n314_n876# 0.41883f
C66 a_n915_7081# AVDD 0.07137f
C67 a_n722_n4252# AVDD 0.91604f
C68 a_n7246_53680# AVDD 19.0667f
C69 a_n2191_3729# MINUS 0.06046f
C70 a_51521_37180# AVDD 19.7915f
C71 a_n314_n876# a_n7496_n2395# 0.06224f
C72 a_n314_n876# AVDD 3.00884f
C73 a_9374_n4648# AVDD 1.224f
C74 m6_n78189_n74849# m7_n78189_n74849# 81.275f
C75 m3_n77751_n74411# m4_n77751_n74411# 0.42115p
C76 a_7669_2986# a_9374_n4648# 0.06823f
C77 a_2417_7081# a_n314_n876# 0.07206f
C78 a_51524_n4820# VOUT 19.1316f
C79 a_n28191_n62820# PLUS 19.1977f
C80 a_n2343_7081# a_n314_n876# 0.07247f
C81 a_n2191_3729# IBIAS 0.38303f
C82 a_n1791_7045# a_n2227_3805# 1.26525f
C83 a_n314_n876# MINUS 0.26316f
C84 a_2893_7081# AVDD 0.069f
C85 a_n2191_3729# m1_n686_n6334# 0.42462f
C86 a_n2191_3729# a_n2227_3805# 1.42728f
C87 a_n1867_7081# AVDD 0.07093f
C88 a_7578_n5569# VOUT 0.33471f
C89 a_51527_n25820# VOUT 19.8298f
C90 m3_n78189_n74849# m4_n78189_n74849# 0.42142p
C91 a_1465_7081# a_n314_n876# 0.07254f
C92 a_n722_n4252# m1_n686_n6334# 0.23704f
C93 a_1623_4206# a_n314_n876# 0.07245f
C94 m5_n77705_n74365# m6_n77609_n74269# 0.17289p
C95 a_n1791_7045# a_n2191_3729# 0.95047f
C96 a_n7496_n2395# VOUT 0.1598f
C97 a_n2227_3805# a_9374_n4648# 0.10225f
C98 a_n2227_3805# a_n314_n876# 1.08527f
C99 a_n7496_n1298# PLUS 0.57722f
C100 AVDD VOUT 3.86948f
C101 a_n2227_3805# a_7669_5842# 0.06914f
C102 a_n65913_n26320# IBIAS 19.5782f
C103 a_n314_276# PLUS 0.2477f
C104 a_1941_7081# AVDD 0.07137f
C105 a_n2811_7081# AVDD 0.06912f
C106 AVDD PLUS 1.96753f
C107 a_n1791_7045# a_9374_n4648# 0.83979f
C108 a_n1791_7045# a_n314_n876# 1.25477f
C109 a_n2191_3729# a_n722_n4252# 0.46935f
C110 a_n49227_53680# MINUS 20.0584f
C111 a_n2191_3729# a_9374_n4648# 0.01919f
C112 m5_n78189_n74849# m6_n78189_n74849# 0.26773p
C113 MINUS PLUS 0.17563f
C114 a_n1791_7045# a_7669_6794# 0.06988f
C115 a_n28215_53180# MINUS 19.1438f
C116 a_13754_53180# AVDD 19.2452f
C117 a_34797_53680# AVDD 19.8224f
C118 a_n2227_3805# VOUT 0.97646f
C119 w_6489_n1941# AVDD 0.04163f
C120 a_n2191_5157# a_n314_276# 0.07207f
C121 PLUS IBIAS 0.0293f
C122 m1_n686_n6334# PLUS 0.02016f
C123 m6_n77609_n74269# m7_n78189_n74849# 52.4849f
C124 a_492_n3852# m1_492_n6334# 0.03122f
C125 a_n2191_3729# VOUT 0.24253f
C126 a_492_n5390# m1_492_n6334# 0.03183f
C127 a_492_n6342# m1_492_n6334# 0.03137f
C128 a_n1791_7045# a_7669_1082# 0.0746f
C129 a_492_n3376# VOUT 0.03213f
C130 m7_n78189_n74849# AVSS 0.20397p
C131 m6_n77609_n74269# AVSS 0.23282p
C132 m6_n78189_n74849# AVSS 0.23435p
C133 m5_n77705_n74365# AVSS 0.17154p
C134 m5_n78189_n74849# AVSS 0.17256p
C135 m4_n77751_n74411# AVSS 0.18129p
C136 m4_n78189_n74849# AVSS 0.18232p
C137 m3_n77751_n74411# AVSS 0.19544p
C138 m3_n78189_n74849# AVSS 0.19654p
C139 m2_n77751_n74411# AVSS 0.21692p
C140 m2_n78189_n74849# AVSS 0.21814p
C141 m1_492_n6334# AVSS 1.42623f
C142 m1_n686_n6334# AVSS 1.40614f
C143 m1_n77751_n74411# AVSS 0.46612p
C144 m1_n78189_n74849# AVSS 0.46765p
C145 a_34774_n62320# AVSS 19.9156f $ **FLOATING
C146 a_13764_n62820# AVSS 19.2666f $ **FLOATING
C147 a_n7223_n62320# AVSS 19.1318f $ **FLOATING
C148 a_51476_n46820# AVSS 19.8731f $ **FLOATING
C149 a_492_n5866# AVSS 0.03034f $ **FLOATING
C150 a_n686_n5866# AVSS 0.03054f $ **FLOATING
C151 a_9374_n4648# AVSS 4.14508f $ **FLOATING
C152 a_7578_n5569# AVSS 4.75877f $ **FLOATING
C153 a_n722_n4252# AVSS 6.6814f $ **FLOATING
C154 a_n7496_n2395# AVSS 6.77414f $ **FLOATING
C155 a_n314_n876# AVSS 3.10706f $ **FLOATING
C156 a_n7496_n1298# AVSS 2.96346f $ **FLOATING
C157 a_n314_276# AVSS 3.82085f $ **FLOATING
C158 a_n2227_3805# AVSS 7.49914f $ **FLOATING
C159 a_n2191_3729# AVSS 15.4068f $ **FLOATING
C160 a_n1791_7045# AVSS 9.81839f $ **FLOATING
.ends
