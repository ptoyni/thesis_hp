* Extracted by KLayout with SG13G2 LVS runset on : 25/06/2025 10:10

.SUBCKT testing_dummies VSS IN VDD
M$1 VSS VSS VDD VSS sg13_lv_nmos L=1u W=4u AS=1.1p AD=0.83p PS=7.1u PD=6.83u
M$2 VDD IN VSS VSS sg13_lv_nmos L=1u W=4u AS=0.76p AD=0.76p PS=4.76u PD=4.76u
.ENDS testing_dummies
