.subckt ota_final VDD VSS
.ends
.end
