.subckt FMD_QNC_ota_final_esd VDD VSS
.ends
.end
