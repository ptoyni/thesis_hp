* Extracted by KLayout with SG13G2 LVS runset on : 25/05/2025 15:29

.SUBCKT sg13g2_buf_1_iso VSS VDD
M$1 VSS \$5 \$1 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.159375p AD=0.247625p
+ PS=1.19u PD=2.29u
M$2 VSS \$1 \$3 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.159375p AD=0.2516p
+ PS=1.19u PD=2.16u
M$3 VDD \$5 \$1 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2051p AD=0.3024p PS=1.52u
+ PD=2.4u
M$4 VDD \$1 \$3 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2051p AD=0.4032p PS=1.52u
+ PD=2.96u
.ENDS sg13g2_buf_1_iso
