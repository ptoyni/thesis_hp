** sch_path: /foss/designs/Thesis/workspace/thesis_hp/Designs/Analog_Inverter/Schematics/Analog_Inverter/testbenches_Analog_Inverter/tb_Analog_Inverter_tran.sch
**.subckt tb_Analog_Inverter_tran
Vdd1 Vdd GND 1.5
Vss1 Vss GND 0
x1 Vdd v_in v_out Vss Analog_Inverter
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt




Vin v_in 0 dc 0 pulse(0 1.5 0 1n 1n 4n 10n)
.control


* Transient analysis
tran 0.01n 20n
save all
let VP=1.5
let per10 = Vp*0.1
let per50 = Vp*0.5
let per90 = Vp*0.9
meas TRAN t_rise  TRIG v(v_out) VAL=per10 rise=2  TARG v(v_out) VAL=per90 rise=2
meas TRAN t_fall  TRIG v(v_out) VAL=per90 fall=2  TARG v(v_out) VAL=per10 fall=2
meas TRAN t_delay  TRIG v(v_in) VAL=per50 rise=1 TARG v(v_out) VAL=per50 fall=1
echo TRAN measurements
print t_delay
print t_rise
print t_fall
echo
*set filetype=binary
*write ./Analog_Inverter/simulations/tb_inv_dc.raw


plot v(v_out) v(v_in)

.endc
.end


**** end user architecture code
**.ends

* expanding   symbol:
*+  /foss/designs/Thesis/workspace/thesis_hp/Designs/Analog_Inverter/Schematics/Analog_Inverter/Analog_Inverter.sym # of pins=4
** sym_path: /foss/designs/Thesis/workspace/thesis_hp/Designs/Analog_Inverter/Schematics/Analog_Inverter/Analog_Inverter.sym
** sch_path: /foss/designs/Thesis/workspace/thesis_hp/Designs/Analog_Inverter/Schematics/Analog_Inverter/Analog_Inverter.sch
.subckt Analog_Inverter vdd vin vout vss
*.ipin vin
*.iopin vdd
*.iopin vss
*.opin vout
XM1 vout vin vdd vdd sg13_lv_pmos w=40u l=0.52u ng=1 m=1
XM2 vout vin vss vss sg13_lv_nmos w=20u l=0.52u ng=1 m=1
.ends

.GLOBAL GND
.end
