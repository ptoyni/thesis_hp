** sch_path: /foss/designs/thesis_hp/designs/otas/1_schematics/foldedcascode_pmos.sch
.SUBCKT foldedcascode_pmos AVDD IBIAS PLUS MINUS VOUT AVSS
*.PININFO PLUS:I MINUS:I AVSS:I IBIAS:I AVDD:I VOUT:O
M1 net6 MINUS net1 AVDD sg13_lv_pmos w=20u l=2u ng=4 m=1
M5 net7 net8 net4 AVSS sg13_lv_nmos w=2u l=2u ng=2 m=1
M2 net4 PLUS net1 AVDD sg13_lv_pmos w=20u l=2u ng=4 m=1
M3 net2 net7 AVDD AVDD sg13_lv_pmos w=13u l=2u ng=2 m=1
M4 net3 net7 AVDD AVDD sg13_lv_pmos w=13u l=2u ng=2 m=1
M7 net7 net9 net2 AVDD sg13_lv_pmos w=8u l=2u ng=4 m=1
M8 VOUT net9 net3 AVDD sg13_lv_pmos w=8u l=2u ng=4 m=1
M6 VOUT net8 net6 AVSS sg13_lv_nmos w=2u l=2u ng=2 m=1
M9 net4 net5 AVSS AVSS sg13_lv_nmos w=4u l=2u ng=2 m=1
M0 net6 net5 AVSS AVSS sg13_lv_nmos w=4u l=2u ng=2 m=1
Mt net1 net10 AVDD AVDD sg13_lv_pmos w=32u l=5u ng=4 m=1
M13 IBIAS net7 net5 AVSS sg13_lv_nmos w=4u l=2u ng=2 m=1
M15 net5 net5 AVSS AVSS sg13_lv_nmos w=4u l=2u ng=1 m=1
M16 net8 net5 AVSS AVSS sg13_lv_nmos w=4u l=2u ng=1 m=1
M14 AVDD net7 net8 AVSS sg13_lv_nmos w=15u l=0.5u ng=2 m=1
M12 net9 net8 AVSS AVSS sg13_lv_nmos w=2u l=2u ng=1 m=1
M10 net9 net9 AVDD AVDD sg13_lv_pmos w=8u l=2u ng=2 m=1
M11 net10 net5 AVSS AVSS sg13_lv_nmos w=4u l=2u ng=1 m=1
Mtb net10 net10 AVDD AVDD sg13_lv_pmos w=28u l=5u ng=4 m=1
M18 net5 AVSS AVSS AVSS sg13_lv_nmos w=4u l=2u ng=1 m=1
M19 AVDD AVSS AVSS AVSS sg13_lv_nmos w=15u l=0.5u ng=2 m=1
M20 net4 AVSS AVSS AVSS sg13_lv_nmos w=4u l=2u ng=2 m=1
M21 net7 AVSS AVSS AVSS sg13_lv_nmos w=2u l=2u ng=2 m=1
M22 VOUT AVSS AVSS AVSS sg13_lv_nmos w=2u l=2u ng=2 m=1
M23 AVDD AVDD net1 AVDD sg13_lv_pmos w=10u l=2u ng=2 m=1
M24 AVDD AVDD net1 AVDD sg13_lv_pmos w=10u l=2u ng=2 m=1
M25 net10 AVSS AVSS AVSS sg13_lv_nmos w=8u l=2u ng=2 m=1
M26 net9 AVSS AVSS AVSS sg13_lv_nmos w=4u l=2u ng=2 m=1
Mtb1 net10 AVDD AVDD AVDD sg13_lv_pmos w=14u l=5u ng=2 m=1
M27 net9 AVDD AVDD AVDD sg13_lv_pmos w=8u l=2u ng=2 m=1
Mt1 AVDD AVDD AVDD AVDD sg13_lv_pmos w=16u l=5u ng=2 m=1
M28 AVDD AVDD AVDD AVDD sg13_lv_pmos w=7.5u l=2u ng=1 m=1
M29 AVDD AVDD AVDD AVDD sg13_lv_pmos w=13u l=2u ng=2 m=1
D3 AVDD AVDD AVSS diodevdd_2kv m=1
D4 AVDD AVDD AVSS diodevss_2kv m=1
D5 AVDD AVSS AVSS diodevdd_2kv m=1
D6 AVDD AVSS AVSS diodevss_2kv m=1
X2 AVSS bondpad
X3 AVDD bondpad
D7 AVDD IBIAS AVSS diodevdd_2kv m=1
D8 AVDD IBIAS AVSS diodevss_2kv m=1
X4 IBIAS bondpad
C2 VOUT AVSS cap_cmim w=25.82e-6 l=25.82e-6 m=1
X1 VOUT bondpad
D1 AVDD VOUT AVSS diodevdd_2kv m=1
D2 AVDD VOUT AVSS diodevss_2kv m=1
X5 PLUS bondpad
X6 MINUS bondpad
D11 AVDD PLUS AVSS diodevdd_2kv m=1
D9 AVDD MINUS AVSS diodevdd_2kv m=1
D12 AVDD PLUS AVSS diodevss_2kv m=1
D10 AVDD MINUS AVSS diodevss_2kv m=1
M30 net8 AVSS AVSS AVSS sg13_lv_nmos w=4u l=2u ng=1 m=1
.ENDS
