* Extracted by KLayout with SG13G2 LVS runset on : 10/07/2025 04:27

.SUBCKT ota_final AVDD IBIAS VOUT MINUS PLUS AVSS
X1 AVDD VOUT \$22047 AVSS sg13_lv_nmos L=0.5u W=15u AS=3.4125p AD=3.4125p
+ PS=20.57u PD=20.57u
X5 AVSS IBIAS IBIAS AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
X9 AVSS IBIAS \$23068 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
X13 AVSS IBIAS \$23067 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
X17 AVSS AVSS \$23210 AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
X18 \$23210 MINUS \$23067 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p
+ PS=6.76u PD=6.76u
X19 \$23067 PLUS \$23491 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p
+ PS=6.76u PD=6.76u
X20 \$23491 AVSS AVSS AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
X25 \$23068 \$22499 \$23069 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
X29 AVSS \$22499 \$23071 AVDD sg13_lv_pmos L=0.5u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
X33 \$21897 VOUT \$22049 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
X35 AVSS AVSS \$21897 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
X36 \$21897 \$21897 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
X37 AVSS \$21897 \$22047 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
X41 AVSS AVSS VOUT AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
X42 VOUT \$22047 \$I560786 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
X45 AVSS AVSS \$I560786 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
X46 \$I560786 \$22499 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
X49 AVSS AVSS \$I560785 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
X50 \$I560785 \$22499 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
X53 AVSS AVSS \$22499 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
X54 \$22499 \$22047 \$I560785 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
X57 AVDD AVDD \$23069 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p
+ PS=11.56u PD=11.56u
X58 \$23069 \$23069 AVDD AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
X59 AVDD \$23069 \$23071 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
X61 AVDD \$23069 \$22049 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
X71 AVDD AVDD \$22499 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p
+ PS=11.56u PD=11.56u
X72 \$22499 \$23071 \$23491 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
X77 AVDD AVDD VOUT AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
X78 VOUT \$23071 \$23210 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
X83 AVDD AVDD \$23210 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
X85 AVDD \$23069 \$23491 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
X87 AVDD \$23069 \$23210 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
.ENDS ota_final
