* NGSPICE file created from complete_schematic_pads_fillers.ext - technology: ihp-sg13g2

.subckt complete_schematic_pads_fillers
X0 a_n7059_10169# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X1 a_981_18638# a_n6059_11418# a_n73946_n58819# a_n73946_n58819# sg13_lv_nmos ad=0.1005p pd=1.34u as=0.1005p ps=1.34u w=0.15u l=10u
X2 vdd a_n7059_10169# a_n7288_16809# vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X3 a_n7289_16017# a_527_15753# rppd l=38.65u w=0.5u
X4 a_n7288_18340# a_528_18033# rppd l=38.65u w=0.71u
X5 a_n73946_n58819# a_5580_15247# a_n7059_10169# a_n73946_n58819# sg13_lv_nmos ad=2.448p pd=15.08u as=1.368p ps=7.58u w=7.2u l=9.75u
X6 a_n6059_10861# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X7 a_n7059_10169# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=3.1875p ps=19.43u w=9.375u l=2.08u
X8 a_4707_16560# vdd vdd vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X9 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X10 vdd a_3822_10479# a_n7059_10169# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X11 vdd a_n7059_10169# a_n7288_16809# vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X12 a_3822_10479# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X13 a_5580_15247# a_3630_15211# a_n73946_n58819# a_n73946_n58819# sg13_lv_nmos ad=0.2448p pd=2.12u as=0.2448p ps=2.12u w=0.72u l=9.75u
X14 vdd a_3822_10479# a_n7059_10169# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X15 vdd a_3822_10479# a_4707_16560# vdd sg13_lv_pmos ad=1.802p pd=11.28u as=1.802p ps=11.28u w=5.3u l=1.95u
X16 a_n73946_n58819# a_n6059_10861# a_n6059_11418# a_n73946_n58819# sg13_lv_nmos ad=0.33915p pd=2.165u as=0.33915p ps=2.165u w=1.785u l=5u
X17 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X18 a_3822_10479# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=3.1875p ps=19.43u w=9.375u l=2.08u
X19 a_4707_16560# vdd vdd vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X20 vdd a_3822_10479# a_n7059_10169# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X21 vdd a_3822_10479# a_3822_10479# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X22 a_n7288_18340# a_n73946_n58819# rppd l=38.65u w=0.71u
X23 vdd a_3822_10479# a_3822_10479# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X24 a_n6059_11418# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X25 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X26 a_n6059_10861# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X27 a_n73946_n58819# a_n7289_16545# a_n7289_16545# a_n73946_n58819# sg13_lv_nmos ad=0.8925p pd=5.93u as=0.49875p ps=3.005u w=2.625u l=5u
X28 a_1804_15931# a_n73946_n58819# cap_cmim l=18.2u w=18.2u
X29 a_n7289_16545# a_n7289_16545# a_n73946_n58819# a_n73946_n58819# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X30 vdd a_3822_10479# a_3822_10479# vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X31 a_n7289_16545# a_n7289_16545# a_n73946_n58819# a_n73946_n58819# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X32 a_n7289_16017# a_527_16281# rppd l=38.65u w=0.5u
X33 vdd a_n7059_10169# a_n6059_10861# vdd sg13_lv_pmos ad=0.6375p pd=4.43u as=0.35625p ps=2.255u w=1.875u l=5u
X34 a_3630_15211# a_n6059_11418# a_4707_16560# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X35 a_n7059_10169# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X36 a_n6059_11418# a_n6059_10861# a_n73946_n58819# a_n73946_n58819# sg13_lv_nmos ad=0.33915p pd=2.165u as=0.33915p ps=2.165u w=1.785u l=5u
X37 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X38 a_n7289_16545# a_n7289_16545# a_n73946_n58819# a_n73946_n58819# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.8925p ps=5.93u w=2.625u l=5u
X39 a_n7288_17727# a_528_18033# rppd l=38.65u w=0.71u
X40 a_n6059_11418# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X41 a_n7288_17115# a_528_16809# rppd l=38.65u w=0.71u
X42 a_n7288_16809# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X43 a_1804_15931# a_981_18638# vdd vdd sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X44 a_5580_15247# a_n6059_10861# a_4707_16560# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X45 a_n7059_10169# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X46 a_n7289_15489# a_527_15753# rppd l=38.65u w=0.5u
X47 a_3822_10479# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X48 vdd a_3822_10479# a_n7059_10169# vdd sg13_lv_pmos ad=3.1875p pd=19.43u as=1.78125p ps=9.755u w=9.375u l=2.08u
X49 vdd a_n7059_10169# a_n6059_11418# vdd sg13_lv_pmos ad=0.6375p pd=4.43u as=0.35625p ps=2.255u w=1.875u l=5u
X50 a_981_18638# a_981_18638# vdd vdd sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X51 a_n7289_15489# a_n6059_10861# rppd l=38.65u w=0.5u
X52 a_n73946_n58819# a_n7289_16545# a_n7289_16545# a_n73946_n58819# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X53 a_3822_10479# a_3822_10479# vdd vdd sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X54 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X55 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X56 vdd a_3822_10479# a_3822_10479# vdd sg13_lv_pmos ad=3.1875p pd=19.43u as=1.78125p ps=9.755u w=9.375u l=2.08u
X57 a_n73946_n58819# a_527_13669# rppd l=38.65u w=3u
X58 a_n7288_16809# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X59 a_n7289_14961# a_n6059_10861# rppd l=38.65u w=0.5u
X60 vdd a_n7059_10169# a_n7288_16809# vdd sg13_lv_pmos ad=0.68p pd=4.68u as=0.38p ps=2.38u w=2u l=5u
X61 a_n6059_11418# a_n6059_10861# a_n73946_n58819# a_n73946_n58819# sg13_lv_nmos ad=0.33915p pd=2.165u as=0.6069p ps=4.25u w=1.785u l=5u
X62 a_n73946_n58819# a_5580_15247# a_n7059_10169# a_n73946_n58819# sg13_lv_nmos ad=1.368p pd=7.58u as=1.368p ps=7.58u w=7.2u l=9.75u
X63 a_n6059_10861# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.6375p ps=4.43u w=1.875u l=5u
X64 a_4707_16560# vdd vdd vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X65 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X66 a_n6059_10861# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X67 a_4707_16560# vdd vdd vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X68 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X69 a_n7059_10169# a_5580_15247# a_n73946_n58819# a_n73946_n58819# sg13_lv_nmos ad=1.368p pd=7.58u as=1.368p ps=7.58u w=7.2u l=9.75u
X70 vdd a_n7059_10169# a_n6059_10861# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X71 a_n6059_11418# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.6375p ps=4.43u w=1.875u l=5u
X72 vdd a_1804_15931# a_n6059_11418# vdd sg13_lv_pmos ad=0.104p pd=1.34u as=0.104p ps=1.34u w=0.2u l=4u
X73 vdd a_981_18638# a_981_18638# vdd sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X74 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X75 a_5580_15247# a_n7059_10169# cap_cmim l=22.29u w=22.29u
X76 a_n6059_11418# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X77 a_5580_15247# a_n6059_10861# a_4707_16560# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X78 vdd a_981_18638# a_1804_15931# vdd sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X79 a_n73946_n58819# a_n7289_16545# a_n7289_16545# a_n73946_n58819# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X80 a_n7288_17115# a_528_17421# rppd l=38.65u w=0.71u
X81 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X82 a_n7289_16545# a_n7289_16545# a_n73946_n58819# a_n73946_n58819# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X83 vdd a_n7059_10169# a_n6059_11418# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X84 vdd a_n7059_10169# a_n6059_10861# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X85 a_n7289_14961# a_527_14697# rppd l=38.65u w=0.5u
X86 vdd vdd a_3630_15211# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X87 a_n73946_n58819# a_n7289_16545# a_n7289_16545# a_n73946_n58819# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X88 a_3630_15211# a_n6059_11418# a_4707_16560# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X89 a_n7288_16809# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.68p ps=4.68u w=2u l=5u
X90 a_n7289_14433# a_527_14697# rppd l=38.65u w=0.5u
X91 vdd a_n7059_10169# a_n6059_10861# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X92 a_n7288_17727# a_528_17421# rppd l=38.65u w=0.71u
X93 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X94 a_n7288_16809# a_n7059_10169# vdd vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X95 vdd vdd a_5580_15247# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X96 a_n7288_16809# a_528_16809# rppd l=38.65u w=0.71u
X97 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X98 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X99 a_n7059_10169# a_5580_15247# a_n73946_n58819# a_n73946_n58819# sg13_lv_nmos ad=1.368p pd=7.58u as=2.448p ps=15.08u w=7.2u l=9.75u
X100 vdd a_n7059_10169# a_n6059_11418# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X101 vdd vdd a_5580_15247# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X102 vdd a_n7059_10169# a_n7288_16809# vdd sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X103 a_n73946_n58819# a_n6059_10861# a_n6059_11418# a_n73946_n58819# sg13_lv_nmos ad=0.6069p pd=4.25u as=0.33915p ps=2.165u w=1.785u l=5u
X104 a_n7289_16545# a_527_16281# rppd l=38.65u w=0.5u
X105 a_n7289_14433# a_527_13669# rppd l=38.65u w=0.5u
X106 a_3630_15211# a_3630_15211# a_n73946_n58819# a_n73946_n58819# sg13_lv_nmos ad=0.2448p pd=2.12u as=0.2448p ps=2.12u w=0.72u l=9.75u
X107 vdd a_n7059_10169# a_n6059_11418# vdd sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X108 vdd vdd a_3630_15211# vdd sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X109 vdd a_n73946_n58819# cap_cmim l=5u w=5u
X110 vdd a_n73946_n58819# cap_cmim l=5u w=5u
C0 a_3822_10479# a_n7059_10169# 3.1169f
C1 a_4707_16560# a_3630_15211# 2.29139f
C2 w_n7489_9836# vdd 0.44088f
C3 a_n7289_16545# a_n6059_11418# 0.4148f
C4 a_n7203_16545# a_527_16281# 0.01946f
C5 w_3320_10081# a_3630_15211# 0.01188f
C6 a_n6059_10861# vdd 7.47803f
C7 a_528_17421# a_n6059_11418# 0.0115f
C8 a_n7202_17115# vdd 0.0101f
C9 a_n7288_16809# a_n7289_14961# 0.01169f
C10 a_n6059_11418# m3_1900_17599# 0.26018f
C11 w_8745_13831# a_5580_15247# 0.01152f
C12 a_n7203_16017# a_n7203_15753# 0.56632f
C13 a_n6059_10861# a_527_15753# 0.02893f
C14 a_n7203_15489# a_n7203_15225# 0.56632f
C15 w_1450_16710# a_n6059_11418# 0.01881f
C16 a_n6059_11418# a_3630_15211# 3.2036f
C17 a_1804_15931# a_5580_15247# 1.05678f
C18 a_n7202_17421# a_n7289_16545# 0.01625f
C19 a_n7202_17115# a_n7202_16809# 0.56632f
C20 a_n6059_10861# a_n7203_15225# 0.03934f
C21 w_3320_16060# a_n6059_10861# 0.0446f
C22 a_528_17421# a_n7202_17421# 0.02797f
C23 a_n7289_16545# a_n7289_16017# 0.02817f
C24 a_n7203_14697# a_n7203_14433# 0.56632f
C25 a_n7288_17727# a_n7202_18033# 0.02797f
C26 a_n7059_10169# vdd 52.2225f
C27 m6_n73506_n58379# m7_n73946_n58819# 49.7261f
C28 a_n7202_18646# a_n7202_18340# 0.56632f
C29 a_n6059_10861# a_5580_15247# 1.86924f
C30 m4_n73648_n58521# m5_n73602_n58475# 0.35175p
C31 a_527_16281# a_527_15753# 0.01716f
C32 a_n7289_16545# a_n7203_16545# 0.52649f
C33 w_1389_15644# a_n6059_11418# 0.01287f
C34 a_3630_15211# a_3822_10479# 0.24066f
C35 m2_n73946_n58819# m3_n73946_n58819# 0.25526p
C36 a_n7203_14961# a_527_14697# 0.01946f
C37 m2_n73648_n58521# m3_n73648_n58521# 0.39679p
C38 w_n7489_9836# a_1804_15931# 0.01251f
C39 a_981_18638# m3_1900_17599# 0.06332f
C40 a_1804_15931# a_n6059_10861# 0.37731f
C41 a_n6059_11418# a_4707_16560# 1.56095f
C42 a_n7289_16545# a_n7203_13669# 1.21239f
C43 a_n7289_15489# a_n7203_15489# 0.01947f
C44 a_528_16809# a_n6059_11418# 0.01664f
C45 a_n7289_16545# vdd 0.36927f
C46 a_n6059_10861# a_n7203_15489# 0.03695f
C47 a_n7289_16017# a_n7203_16017# 0.01946f
C48 a_n7289_16545# a_n7203_14961# 0.05896f
C49 w_1450_16710# a_981_18638# 0.01837f
C50 a_5580_15247# a_n7059_10169# 29.8065f
C51 a_527_14697# a_527_13669# 0.01716f
C52 a_n7202_18340# a_n7202_18033# 0.5628f
C53 m3_1900_17599# vdd 0.09726f
C54 w_n7489_9836# a_n6059_10861# 0.01778f
C55 a_n7202_18646# vdd 0.05279f
C56 a_n7289_16545# a_527_15753# 0.01099f
C57 a_n7202_16809# a_n7289_16545# 0.11069f
C58 w_1450_16710# vdd 0.13817f
C59 a_3630_15211# vdd 4.89658f
C60 a_n7289_16545# a_527_13669# 0.01975f
C61 a_4707_16560# a_3822_10479# 1.1372f
C62 a_n7202_17727# a_n7289_16545# 0.04457f
C63 a_n7288_17115# a_n7288_16809# 0.0308f
C64 a_n7289_16545# a_n7203_15225# 0.25983f
C65 a_n7202_17727# a_528_17421# 0.02797f
C66 w_3320_10081# a_3822_10479# 0.04216f
C67 a_1804_15931# a_n7059_10169# 0.27209f
C68 a_n7288_18340# a_n7202_18646# 0.02797f
C69 a_n7288_16809# a_n7203_13669# 0.02294f
C70 m3_n73946_n58819# m4_n73946_n58819# 0.25526p
C71 w_n7489_9836# a_n7059_10169# 0.07536f
C72 a_n7203_14433# a_n7203_13669# 0.56632f
C73 a_n7288_16809# vdd 5.7108f
C74 w_1389_15644# vdd 0.08151f
C75 a_n6059_10861# a_n7059_10169# 2.09172f
C76 m3_n73648_n58521# m4_n73648_n58521# 0.39679p
C77 w_3320_16060# a_3630_15211# 0.05123f
C78 a_527_16281# a_n7203_16281# 0.01946f
C79 a_n7202_18033# vdd 0.02044f
C80 a_n7288_17727# a_n7288_17115# 0.01716f
C81 a_n7289_14961# a_n7203_14961# 0.01946f
C82 a_n7203_16017# a_527_15753# 0.01946f
C83 a_5580_15247# a_3630_15211# 2.48082f
C84 a_n7288_16809# a_n7202_16809# 0.05671f
C85 a_n7289_16545# a_1804_15931# 0.05182f
C86 a_4707_16560# vdd 2.39323f
C87 a_n6059_10861# a_527_14697# 0.0297f
C88 a_n7203_14433# a_527_13669# 0.01946f
C89 a_n7289_16545# a_n7203_15489# 0.07779f
C90 a_n7202_18033# a_n7202_17727# 0.56632f
C91 w_3320_10081# vdd 0.29549f
C92 a_1804_15931# m3_1900_17599# 0.19258f
C93 a_981_18638# a_n6059_11418# 0.36328f
C94 a_n7203_14961# a_n7203_14697# 0.56632f
C95 a_527_15753# a_n7203_15753# 0.01946f
C96 w_n7489_9836# a_n7289_16545# 0.04233f
C97 a_n7289_14961# a_n7203_15225# 0.01946f
C98 w_1450_16710# a_1804_15931# 0.02595f
C99 a_n7289_16545# a_n6059_10861# 0.08938f
C100 a_n6059_11418# a_n7203_13669# 0.01352f
C101 a_n7202_17115# a_n7289_16545# 0.14683f
C102 a_528_16809# a_n7202_16809# 0.02797f
C103 a_n6059_10861# m3_1900_17599# 0.01692f
C104 a_n6059_11418# vdd 6.42134f
C105 w_3320_16060# a_4707_16560# 0.02689f
C106 a_n7288_17115# a_n7202_17421# 0.02797f
C107 a_n7289_16545# a_n7203_16281# 0.12328f
C108 a_n7288_17727# a_n7202_17727# 0.02797f
C109 a_528_18033# a_528_17421# 0.01716f
C110 a_981_18638# a_n7202_18340# 0.0122f
C111 a_n7288_18340# a_n7288_17727# 0.01705f
C112 a_n6059_10861# a_3630_15211# 2.14089f
C113 a_4707_16560# a_5580_15247# 1.867f
C114 a_n6059_11418# a_527_15753# 0.01654f
C115 a_n7289_16545# a_527_16281# 0.03485f
C116 a_n7202_16809# a_n6059_11418# 0.01976f
C117 w_1389_15644# a_1804_15931# 0.03719f
C118 w_3320_10081# a_5580_15247# 0.01392f
C119 a_n7289_16545# a_n7059_10169# 0.14068f
C120 w_3320_16060# a_n6059_11418# 0.01719f
C121 a_3822_10479# vdd 55.6035f
C122 a_n7202_18340# vdd 0.1303f
C123 a_n7288_16809# a_n7289_15489# 0.01114f
C124 w_n7489_9836# a_n7288_16809# 0.02439f
C125 a_n7288_16809# a_n6059_10861# 1.54398f
C126 w_1389_15644# a_n6059_10861# 0.02246f
C127 m1_n73946_n58819# m2_n73946_n58819# 0.25526p
C128 a_n6059_11418# a_5580_15247# 0.6702f
C129 a_n7289_15489# a_n7289_14961# 0.01718f
C130 a_n7203_15753# a_n7203_15489# 0.56632f
C131 m1_n73648_n58521# m2_n73648_n58521# 0.39679p
C132 a_n7288_16809# a_n7289_14433# 0.01186f
C133 a_n7203_16281# a_n7203_16017# 0.56632f
C134 a_n7202_17727# a_n7202_17421# 0.56632f
C135 a_n7289_15489# a_n7203_15753# 0.01947f
C136 a_n7289_14433# a_n7203_14433# 0.01946f
C137 a_528_18033# a_n7202_18033# 0.02797f
C138 m6_n73946_n58819# m7_n73946_n58819# 49.2286f
C139 a_n7289_14961# a_n7289_14433# 0.01716f
C140 a_981_18638# vdd 2.62737f
C141 a_n7288_18340# a_n7202_18340# 0.02797f
C142 m4_n73946_n58819# m5_n73946_n58819# 0.25526p
C143 a_n6059_10861# a_4707_16560# 1.00293f
C144 a_n7202_16809# a_n7203_16545# 0.56625f
C145 w_3320_10081# a_n6059_10861# 0.02816f
C146 a_n6059_11418# a_1804_15931# 0.92177f
C147 a_5580_15247# a_3822_10479# 0.94919f
C148 a_n7202_17115# a_528_16809# 0.02797f
C149 a_n7203_13669# vdd 0.02433f
C150 a_n7288_16809# a_n7059_10169# 9.48469f
C151 a_n7289_14433# a_n7203_14697# 0.01946f
C152 m5_n73602_n58475# m6_n73506_n58379# 0.1638p
C153 w_n7489_9836# a_n6059_11418# 0.04419f
C154 w_8745_13831# a_3822_10479# 0.03192f
C155 a_n6059_11418# a_n6059_10861# 7.74189f
C156 a_527_15753# vdd 0.01523f
C157 a_528_16809# a_527_16281# 0.01695f
C158 a_527_13669# a_n7203_13669# 0.12082f
C159 a_528_18033# a_n6059_11418# 0.01068f
C160 a_n7202_17727# vdd 0.0889f
C161 w_3320_10081# a_n7059_10169# 0.02273f
C162 a_n7203_15225# a_n7203_14961# 0.56632f
C163 w_3320_16060# vdd 0.93984f
C164 a_n7289_16545# a_n7203_16017# 0.08032f
C165 a_n7288_16809# a_n7289_16545# 0.6914f
C166 a_n7289_16017# a_n7289_15489# 0.01718f
C167 a_5580_15247# vdd 10.2641f
C168 a_n6059_10861# a_3822_10479# 0.13837f
C169 a_n7289_16545# a_n7203_14433# 0.18378f
C170 a_n7202_17421# a_n7202_17115# 0.56632f
C171 a_n6059_11418# a_n7059_10169# 1.861f
C172 a_981_18638# a_1804_15931# 1.48658f
C173 a_527_14697# a_n7203_14697# 0.01946f
C174 a_n7202_18340# a_528_18033# 0.02797f
C175 m5_n73946_n58819# m6_n73946_n58819# 0.16216p
C176 a_n7289_16545# a_n7203_15753# 0.28841f
C177 a_n7289_16017# a_n7203_16281# 0.01946f
C178 w_8745_13831# vdd 0.12012f
C179 a_1804_15931# vdd 4.9863f
C180 a_n7289_16545# a_n7203_14697# 0.10236f
C181 w_3320_16060# a_5580_15247# 0.1037f
C182 a_n7288_17115# a_n7202_17115# 0.02797f
C183 a_528_17421# a_528_16809# 0.01716f
C184 a_981_18638# a_n6059_10861# 0.01619f
C185 a_n7203_16545# a_n7203_16281# 0.56632f
C186 m7_n73946_n58819# a_n73946_n58819# 0.19004p
C187 m6_n73506_n58379# a_n73946_n58819# 0.21706p
C188 m6_n73946_n58819# a_n73946_n58819# 0.21838p
C189 m5_n73602_n58475# a_n73946_n58819# 0.15994p
C190 m5_n73946_n58819# a_n73946_n58819# 0.1608p
C191 m4_n73648_n58521# a_n73946_n58819# 0.16903p
C192 m4_n73946_n58819# a_n73946_n58819# 0.16989p
C193 m3_1900_17599# a_n73946_n58819# 0.07675f
C194 m3_n73648_n58521# a_n73946_n58819# 0.18222p
C195 m3_n73946_n58819# a_n73946_n58819# 0.18315p
C196 m2_n73648_n58521# a_n73946_n58819# 0.20225p
C197 m2_n73946_n58819# a_n73946_n58819# 0.20328p
C198 m1_n73648_n58521# a_n73946_n58819# 0.43674p
C199 m1_n73946_n58819# a_n73946_n58819# 0.36419p
C200 a_n7059_10169# a_n73946_n58819# 8.38806f $ **FLOATING
C201 a_n7203_13669# a_n73946_n58819# 13.2658f
C202 a_527_13669# a_n73946_n58819# 0.57903f $ **FLOATING
C203 a_n7203_14433# a_n73946_n58819# 3.81224f
C204 a_n7203_14697# a_n73946_n58819# 3.80717f
C205 a_n7289_14433# a_n73946_n58819# 0.26883f $ **FLOATING
C206 a_527_14697# a_n73946_n58819# 0.25188f $ **FLOATING
C207 a_n7203_14961# a_n73946_n58819# 3.80196f
C208 a_n7203_15225# a_n73946_n58819# 3.79878f
C209 a_n7289_14961# a_n73946_n58819# 0.25151f $ **FLOATING
C210 a_n7203_15489# a_n73946_n58819# 3.79878f
C211 a_n7203_15753# a_n73946_n58819# 3.79878f
C212 a_n7289_15489# a_n73946_n58819# 0.25183f $ **FLOATING
C213 a_527_15753# a_n73946_n58819# 0.23297f $ **FLOATING
C214 a_n7203_16017# a_n73946_n58819# 3.79842f
C215 a_n7203_16281# a_n73946_n58819# 3.79851f
C216 a_n7289_16017# a_n73946_n58819# 0.25103f $ **FLOATING
C217 a_3630_15211# a_n73946_n58819# 6.88509f $ **FLOATING
C218 a_5580_15247# a_n73946_n58819# 45.1225f $ **FLOATING
C219 a_4707_16560# a_n73946_n58819# 2.37087f $ **FLOATING
C220 a_n6059_10861# a_n73946_n58819# 15.2842f $ **FLOATING
C221 a_1804_15931# a_n73946_n58819# 16.217f $ **FLOATING
C222 a_n6059_11418# a_n73946_n58819# 10.3529f $ **FLOATING
C223 a_527_16281# a_n73946_n58819# 0.28604f $ **FLOATING
C224 a_n7203_16545# a_n73946_n58819# 3.79788f
C225 a_n7289_16545# a_n73946_n58819# 37.5098f $ **FLOATING
C226 a_n7202_16809# a_n73946_n58819# 4.50777f
C227 a_528_16809# a_n73946_n58819# 0.34584f $ **FLOATING
C228 a_n7202_17115# a_n73946_n58819# 4.50921f
C229 a_n7202_17421# a_n73946_n58819# 4.50869f
C230 a_n7288_17115# a_n73946_n58819# 0.30345f $ **FLOATING
C231 a_528_17421# a_n73946_n58819# 0.34565f $ **FLOATING
C232 a_n7202_17727# a_n73946_n58819# 4.50921f
C233 a_n7202_18033# a_n73946_n58819# 4.51531f
C234 a_n7288_17727# a_n73946_n58819# 0.30405f $ **FLOATING
C235 a_528_18033# a_n73946_n58819# 0.36381f $ **FLOATING
C236 a_n7202_18340# a_n73946_n58819# 4.55105f
C237 a_981_18638# a_n73946_n58819# 1.18638f $ **FLOATING
C238 a_n7202_18646# a_n73946_n58819# 5.24632f
C239 a_n7288_18340# a_n73946_n58819# 0.3202f $ **FLOATING
C240 w_n7489_9836# a_n73946_n58819# 0.2142f
C241 w_3320_10081# a_n73946_n58819# 0.10287f
C242 w_8745_13831# a_n73946_n58819# 0.02418f
C243 w_3320_16060# a_n73946_n58819# 0.11949f
C244 w_1450_16710# a_n73946_n58819# 0.03111f
.ends
