* NGSPICE file created from full_bandgap.ext - technology: ihp-sg13g2

.subckt full_bandgap vss VBG vdd iout
X0 a_n7059_10169# a_3822_10479# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X1 a_981_18638# a_n6059_11418# a_n74040_n58072# a_n74040_n58072# sg13_lv_nmos ad=0.1005p pd=1.34u as=0.1005p ps=1.34u w=0.15u l=10u
X2 dw_n7489_9836# a_n7059_10169# a_n7288_16809# dw_n7489_9836# sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X3 a_n7289_16017# a_527_15753# rppd l=38.65u w=0.5u
X4 a_n7288_18340# a_528_18033# rppd l=38.65u w=0.71u
X5 a_n74040_n58072# a_5580_15247# a_n7059_10169# a_n74040_n58072# sg13_lv_nmos ad=2.448p pd=15.08u as=1.368p ps=7.58u w=7.2u l=9.75u
X6 a_n6059_10861# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X7 a_n7059_10169# a_3822_10479# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=3.1875p ps=19.43u w=9.375u l=2.08u
X8 a_4707_16560# dw_n7489_9836# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X9 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X10 dw_n7489_9836# a_3822_10479# a_n7059_10169# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X11 dw_n7489_9836# a_n7059_10169# a_n7288_16809# dw_n7489_9836# sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X12 a_3822_10479# a_3822_10479# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X13 a_5580_15247# a_3630_15211# a_n74040_n58072# a_n74040_n58072# sg13_lv_nmos ad=0.2448p pd=2.12u as=0.2448p ps=2.12u w=0.72u l=9.75u
X14 dw_n7489_9836# a_3822_10479# a_n7059_10169# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X15 dw_n7489_9836# a_3822_10479# a_4707_16560# dw_n7489_9836# sg13_lv_pmos ad=1.802p pd=11.28u as=1.802p ps=11.28u w=5.3u l=1.95u
X16 a_n74040_n58072# a_n6059_10861# a_n6059_11418# a_n74040_n58072# sg13_lv_nmos ad=0.33915p pd=2.165u as=0.33915p ps=2.165u w=1.785u l=5u
X17 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X18 a_3822_10479# a_3822_10479# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=3.1875p ps=19.43u w=9.375u l=2.08u
X19 a_4707_16560# dw_n7489_9836# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X20 dw_n7489_9836# a_3822_10479# a_n7059_10169# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X21 dw_n7489_9836# a_3822_10479# a_3822_10479# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X22 a_n7288_18340# a_n74040_n58072# rppd l=38.65u w=0.71u
X23 dw_n7489_9836# a_3822_10479# a_3822_10479# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X24 a_n6059_11418# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X25 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X26 a_n6059_10861# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X27 a_n74040_n58072# a_n7289_16545# a_n7289_16545# a_n74040_n58072# sg13_lv_nmos ad=0.8925p pd=5.93u as=0.49875p ps=3.005u w=2.625u l=5u
X28 a_1804_15931# a_n74040_n58072# cap_cmim l=18.2u w=18.2u
X29 a_n7289_16545# a_n7289_16545# a_n74040_n58072# a_n74040_n58072# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X30 dw_n7489_9836# a_3822_10479# a_3822_10479# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X31 a_n7289_16545# a_n7289_16545# a_n74040_n58072# a_n74040_n58072# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X32 a_n7289_16017# a_527_16281# rppd l=38.65u w=0.5u
X33 dw_n7489_9836# a_n7059_10169# a_n6059_10861# dw_n7489_9836# sg13_lv_pmos ad=0.6375p pd=4.43u as=0.35625p ps=2.255u w=1.875u l=5u
X34 a_3630_15211# a_n6059_11418# a_4707_16560# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X35 a_n7059_10169# a_3822_10479# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X36 a_n6059_11418# a_n6059_10861# a_n74040_n58072# a_n74040_n58072# sg13_lv_nmos ad=0.33915p pd=2.165u as=0.33915p ps=2.165u w=1.785u l=5u
X37 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X38 a_n7289_16545# a_n7289_16545# a_n74040_n58072# a_n74040_n58072# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.8925p ps=5.93u w=2.625u l=5u
X39 a_n7288_17727# a_528_18033# rppd l=38.65u w=0.71u
X40 a_n6059_11418# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X41 a_n7288_17115# a_528_16809# rppd l=38.65u w=0.71u
X42 a_n7288_16809# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X43 a_1804_15931# a_981_18638# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X44 a_5580_15247# a_n6059_10861# a_4707_16560# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X45 a_n7059_10169# a_3822_10479# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X46 a_n7289_15489# a_527_15753# rppd l=38.65u w=0.5u
X47 a_3822_10479# a_3822_10479# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X48 dw_n7489_9836# a_3822_10479# a_n7059_10169# dw_n7489_9836# sg13_lv_pmos ad=3.1875p pd=19.43u as=1.78125p ps=9.755u w=9.375u l=2.08u
X49 dw_n7489_9836# a_n7059_10169# a_n6059_11418# dw_n7489_9836# sg13_lv_pmos ad=0.6375p pd=4.43u as=0.35625p ps=2.255u w=1.875u l=5u
X50 a_981_18638# a_981_18638# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X51 a_n7289_15489# a_n6059_10861# rppd l=38.65u w=0.5u
X52 a_n74040_n58072# a_n7289_16545# a_n7289_16545# a_n74040_n58072# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X53 a_3822_10479# a_3822_10479# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.78125p pd=9.755u as=1.78125p ps=9.755u w=9.375u l=2.08u
X54 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X55 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X56 dw_n7489_9836# a_3822_10479# a_3822_10479# dw_n7489_9836# sg13_lv_pmos ad=3.1875p pd=19.43u as=1.78125p ps=9.755u w=9.375u l=2.08u
X57 a_n74040_n58072# a_527_13669# rppd l=38.65u w=3u
X58 a_n7288_16809# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X59 a_n7289_14961# a_n6059_10861# rppd l=38.65u w=0.5u
X60 dw_n7489_9836# a_n7059_10169# a_n7288_16809# dw_n7489_9836# sg13_lv_pmos ad=0.68p pd=4.68u as=0.38p ps=2.38u w=2u l=5u
X61 a_n6059_11418# a_n6059_10861# a_n74040_n58072# a_n74040_n58072# sg13_lv_nmos ad=0.33915p pd=2.165u as=0.6069p ps=4.25u w=1.785u l=5u
X62 a_n74040_n58072# a_5580_15247# a_n7059_10169# a_n74040_n58072# sg13_lv_nmos ad=1.368p pd=7.58u as=1.368p ps=7.58u w=7.2u l=9.75u
X63 a_n6059_10861# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.6375p ps=4.43u w=1.875u l=5u
X64 a_4707_16560# dw_n7489_9836# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X65 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X66 a_n6059_10861# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X67 a_4707_16560# dw_n7489_9836# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X68 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X69 a_n7059_10169# a_5580_15247# a_n74040_n58072# a_n74040_n58072# sg13_lv_nmos ad=1.368p pd=7.58u as=1.368p ps=7.58u w=7.2u l=9.75u
X70 dw_n7489_9836# a_n7059_10169# a_n6059_10861# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X71 a_n6059_11418# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.6375p ps=4.43u w=1.875u l=5u
X72 dw_n7489_9836# a_1804_15931# a_n6059_11418# dw_n7489_9836# sg13_lv_pmos ad=0.104p pd=1.34u as=0.104p ps=1.34u w=0.2u l=4u
X73 dw_n7489_9836# a_981_18638# a_981_18638# dw_n7489_9836# sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X74 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X75 a_5580_15247# a_n7059_10169# cap_cmim l=22.29u w=22.29u
X76 a_n6059_11418# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X77 a_5580_15247# a_n6059_10861# a_4707_16560# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X78 dw_n7489_9836# a_981_18638# a_1804_15931# dw_n7489_9836# sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=1u
X79 a_n74040_n58072# a_n7289_16545# a_n7289_16545# a_n74040_n58072# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X80 a_n7288_17115# a_528_17421# rppd l=38.65u w=0.71u
X81 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X82 a_n7289_16545# a_n7289_16545# a_n74040_n58072# a_n74040_n58072# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X83 dw_n7489_9836# a_n7059_10169# a_n6059_11418# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X84 dw_n7489_9836# a_n7059_10169# a_n6059_10861# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X85 a_n7289_14961# a_527_14697# rppd l=38.65u w=0.5u
X86 dw_n7489_9836# dw_n7489_9836# a_3630_15211# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X87 a_n74040_n58072# a_n7289_16545# a_n7289_16545# a_n74040_n58072# sg13_lv_nmos ad=0.49875p pd=3.005u as=0.49875p ps=3.005u w=2.625u l=5u
X88 a_3630_15211# a_n6059_11418# a_4707_16560# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X89 a_n7288_16809# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.38p pd=2.38u as=0.68p ps=4.68u w=2u l=5u
X90 a_n7289_14433# a_527_14697# rppd l=38.65u w=0.5u
X91 dw_n7489_9836# a_n7059_10169# a_n6059_10861# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X92 a_n7288_17727# a_528_17421# rppd l=38.65u w=0.71u
X93 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X94 a_n7288_16809# a_n7059_10169# dw_n7489_9836# dw_n7489_9836# sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X95 dw_n7489_9836# dw_n7489_9836# a_5580_15247# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X96 a_n7288_16809# a_528_16809# rppd l=38.65u w=0.71u
X97 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X98 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X99 a_n7059_10169# a_5580_15247# a_n74040_n58072# a_n74040_n58072# sg13_lv_nmos ad=1.368p pd=7.58u as=2.448p ps=15.08u w=7.2u l=9.75u
X100 dw_n7489_9836# a_n7059_10169# a_n6059_11418# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X101 dw_n7489_9836# dw_n7489_9836# a_5580_15247# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X102 dw_n7489_9836# a_n7059_10169# a_n7288_16809# dw_n7489_9836# sg13_lv_pmos ad=0.38p pd=2.38u as=0.38p ps=2.38u w=2u l=5u
X103 a_n74040_n58072# a_n6059_10861# a_n6059_11418# a_n74040_n58072# sg13_lv_nmos ad=0.6069p pd=4.25u as=0.33915p ps=2.165u w=1.785u l=5u
X104 a_n7289_16545# a_527_16281# rppd l=38.65u w=0.5u
X105 a_n7289_14433# a_527_13669# rppd l=38.65u w=0.5u
X106 a_3630_15211# a_3630_15211# a_n74040_n58072# a_n74040_n58072# sg13_lv_nmos ad=0.2448p pd=2.12u as=0.2448p ps=2.12u w=0.72u l=9.75u
X107 dw_n7489_9836# a_n7059_10169# a_n6059_11418# dw_n7489_9836# sg13_lv_pmos ad=0.35625p pd=2.255u as=0.35625p ps=2.255u w=1.875u l=5u
X108 dw_n7489_9836# dw_n7489_9836# a_3630_15211# dw_n7489_9836# sg13_lv_pmos ad=1.2376p pd=7.96u as=1.2376p ps=7.96u w=3.64u l=3.7u
X109 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
X110 dw_n7489_9836# a_n74040_n58072# cap_cmim l=5u w=5u
C0 a_n7203_14433# a_n7289_14433# 0.01946f
C1 a_n7203_14961# a_n7289_16545# 0.25927f
C2 a_527_15753# a_n7289_16545# 0.01192f
C3 a_n7202_17421# a_n7202_17727# 0.56632f
C4 a_n7289_16545# a_n7203_16281# 0.46335f
C5 a_3822_10479# a_n7059_10169# 3.85873f
C6 a_528_17421# a_528_16809# 0.01716f
C7 a_n7203_14433# a_n7203_13669# 0.56632f
C8 a_n6059_11418# a_n7289_16545# 0.66075f
C9 a_n7203_14433# a_n7203_14697# 0.56632f
C10 a_528_18033# a_n7202_18033# 0.02797f
C11 a_n7202_16809# a_n7203_16545# 0.56625f
C12 w_n7489_9836# a_n6059_11418# 0.04419f
C13 dw_n7489_9836# a_n7202_18340# 0.1303f
C14 m4_n74040_n58072# m3_n74040_n58072# 0.39453p
C15 dw_n7489_9836# a_527_15753# 0.01523f
C16 a_3630_15211# a_n6059_10861# 2.21895f
C17 w_3320_10081# a_n7059_10169# 0.03712f
C18 dw_n7489_9836# a_n6059_11418# 6.81155f
C19 w_1450_16710# a_1804_15931# 0.02886f
C20 a_5580_15247# a_n7059_10169# 32.0404f
C21 w_8745_13831# a_4707_16560# 0.01171f
C22 m2_n74040_n58072# m1_n74040_n58072# 0.39453p
C23 dw_n7489_9836# a_3630_15211# 5.91142f
C24 a_n6059_11418# a_1804_15931# 1.06328f
C25 a_n7289_16017# a_n7289_15489# 0.01718f
C26 a_n7203_15489# a_n7203_15225# 0.56632f
C27 a_n7203_15489# a_n7203_15753# 0.56632f
C28 a_n7202_18033# a_n7288_17727# 0.02797f
C29 a_n7289_14433# a_n7203_14697# 0.01946f
C30 a_n7202_17115# a_n7202_16809# 0.56632f
C31 a_3822_10479# w_3320_10081# 0.06138f
C32 a_527_16281# a_n7289_16545# 0.03573f
C33 a_3822_10479# a_5580_15247# 1.0066f
C34 m3_n73602_n57634# m2_n73602_n57634# 0.39413p
C35 a_n6059_11418# a_528_16809# 0.02012f
C36 a_527_14697# a_n7203_14697# 0.01946f
C37 a_n7203_15489# a_n6059_10861# 0.03922f
C38 a_n6059_11418# m3_1900_17599# 0.26018f
C39 w_3320_10081# a_5580_15247# 0.01939f
C40 a_n7203_15489# a_n7289_16545# 0.27748f
C41 w_8745_13831# dw_n7489_9836# 0.12231f
C42 a_n7202_17727# a_n7289_16545# 0.04493f
C43 a_n6059_11418# a_528_17421# 0.01278f
C44 a_n7202_18646# dw_n7489_9836# 0.19793f
C45 a_n7202_17421# a_n7202_17115# 0.56632f
C46 dw_n7489_9836# a_n7202_17727# 0.0906f
C47 a_n6059_11418# a_n7203_13669# 0.02588f
C48 a_n7203_14697# a_n7203_14961# 0.56632f
C49 a_5580_15247# w_3320_16060# 0.12191f
C50 a_527_14697# a_n7203_14961# 0.01946f
C51 a_n7059_10169# a_n6059_10861# 3.10863f
C52 a_n7289_14961# a_n7289_15489# 0.01718f
C53 a_527_15753# a_n7203_16017# 0.01946f
C54 m6_n73460_n57492# m5_n73556_n57588# 0.16179p
C55 a_n7203_16017# a_n7203_16281# 0.56632f
C56 a_n7288_18340# a_n7202_18340# 0.02797f
C57 a_n6059_11418# a_n7203_16017# 0.01623f
C58 m6_n73460_n57492# m7_n74040_n58072# 49.114f
C59 a_n7059_10169# a_n7289_16545# 0.19248f
C60 a_3822_10479# a_4707_16560# 1.21741f
C61 w_n7489_9836# a_n7059_10169# 0.0763f
C62 a_527_16281# a_528_16809# 0.01695f
C63 w_1450_16710# a_n6059_11418# 0.02162f
C64 dw_n7489_9836# a_n7059_10169# 53.6649f
C65 a_527_13669# a_n7289_16545# 0.0393f
C66 a_5580_15247# a_4707_16560# 2.20926f
C67 a_n7289_16545# a_n7203_16545# 0.57323f
C68 a_n7289_16017# a_n7289_16545# 0.03605f
C69 a_n7289_15489# a_n7203_15753# 0.01947f
C70 a_527_15753# a_n6059_11418# 0.01738f
C71 a_n7202_16809# a_n7289_16545# 0.31907f
C72 a_3822_10479# a_n6059_10861# 0.1504f
C73 a_n7059_10169# a_1804_15931# 0.35354f
C74 a_981_18638# a_n6059_10861# 0.01705f
C75 a_n7059_10169# a_n7288_16809# 10.5491f
C76 a_n7289_16545# a_n7202_18033# 0.02918f
C77 dw_n7489_9836# a_n7202_16809# 0.01247f
C78 m4_n74040_n58072# m5_n74040_n58072# 0.39453p
C79 a_4707_16560# w_3320_16060# 0.05243f
C80 a_528_17421# a_n7202_17727# 0.02797f
C81 w_3320_10081# a_n6059_10861# 0.03529f
C82 m6_n74040_n58072# m7_n74040_n58072# 76.089f
C83 a_5580_15247# a_n6059_10861# 1.95475f
C84 a_n6059_11418# a_3630_15211# 3.28258f
C85 m3_n73602_n57634# m4_n73602_n57634# 0.39413p
C86 a_3822_10479# dw_n7489_9836# 57.1203f
C87 dw_n7489_9836# a_n7202_18033# 0.10885f
C88 dw_n7489_9836# a_981_18638# 2.65435f
C89 a_n7289_15489# a_n7289_16545# 0.01143f
C90 a_n7203_15225# a_n7289_14961# 0.01946f
C91 dw_n7489_9836# a_n7288_17727# 0.01227f
C92 a_n7288_16809# a_n7289_16017# 0.02643f
C93 a_n7202_17115# a_n7289_16545# 0.14683f
C94 a_527_13669# a_n7203_14433# 0.01946f
C95 a_n7202_16809# a_n7288_16809# 0.06913f
C96 w_3320_10081# dw_n7489_9836# 0.29549f
C97 dw_n7489_9836# a_5580_15247# 11.6825f
C98 a_n7202_17421# a_n7289_16545# 0.07627f
C99 dw_n7489_9836# a_n7202_17115# 0.01249f
C100 w_3320_16060# a_n6059_10861# 0.06145f
C101 a_n7202_18646# a_n7288_18340# 0.02797f
C102 a_981_18638# a_1804_15931# 1.49127f
C103 a_527_15753# a_527_16281# 0.01716f
C104 a_n7202_17421# dw_n7489_9836# 0.01249f
C105 a_527_16281# a_n7203_16281# 0.01946f
C106 a_528_17421# a_528_18033# 0.01716f
C107 a_n7289_14961# a_n7289_16545# 0.01076f
C108 a_n7202_16809# a_528_16809# 0.02797f
C109 a_5580_15247# a_1804_15931# 1.05678f
C110 a_n7288_16809# a_n7289_15489# 0.02618f
C111 w_1389_15644# a_n6059_10861# 0.0227f
C112 dw_n7489_9836# w_3320_16060# 0.9738f
C113 a_n7202_18646# a_n7202_18340# 0.56632f
C114 a_n7288_17115# a_n7288_17727# 0.01716f
C115 a_4707_16560# a_n6059_10861# 1.04184f
C116 a_981_18638# m3_1900_17599# 0.06332f
C117 a_527_13669# a_n7203_13669# 0.12082f
C118 a_n7203_15225# a_n6059_10861# 0.03934f
C119 w_1389_15644# dw_n7489_9836# 0.08151f
C120 a_n7202_17115# a_n7288_17115# 0.02797f
C121 a_527_14697# a_527_13669# 0.01716f
C122 a_n7203_15225# a_n7289_16545# 0.26585f
C123 a_n7289_16545# a_n7203_15753# 0.3003f
C124 a_n7202_17115# a_528_16809# 0.02797f
C125 dw_n7489_9836# a_4707_16560# 3.4745f
C126 a_n7289_14961# a_n7288_16809# 0.01836f
C127 a_n7202_17421# a_n7288_17115# 0.02797f
C128 a_n7203_16017# a_n7289_16017# 0.01946f
C129 a_n6059_11418# a_n7059_10169# 2.78705f
C130 w_1389_15644# a_1804_15931# 0.04245f
C131 a_n7202_18340# a_528_18033# 0.02797f
C132 a_n7289_16545# a_n6059_10861# 0.0901f
C133 a_n6059_11418# a_528_18033# 0.01068f
C134 a_n7202_17421# a_528_17421# 0.02797f
C135 w_n7489_9836# a_n6059_10861# 0.01847f
C136 a_n6059_11418# a_527_13669# 0.01087f
C137 dw_n7489_9836# a_n6059_10861# 8.03346f
C138 a_n7203_16281# a_n7203_16545# 0.56632f
C139 w_n7489_9836# a_n7289_16545# 0.04233f
C140 a_n7288_18340# a_n7288_17727# 0.01705f
C141 w_1450_16710# a_981_18638# 0.01837f
C142 a_n7289_16017# a_n7203_16281# 0.01946f
C143 dw_n7489_9836# a_n7289_16545# 0.4447f
C144 a_n6059_11418# a_n7202_16809# 0.03367f
C145 w_n7489_9836# dw_n7489_9836# 0.44118f
C146 a_n7202_18340# a_n7202_18033# 0.5628f
C147 a_1804_15931# a_n6059_10861# 0.63328f
C148 a_n7289_14961# a_n7289_14433# 0.01716f
C149 a_n7202_18340# a_981_18638# 0.0122f
C150 a_n7288_16809# a_n6059_10861# 1.54398f
C151 a_n6059_11418# a_981_18638# 0.36385f
C152 a_1804_15931# a_n7289_16545# 0.07823f
C153 a_n7288_16809# a_n7289_16545# 0.71412f
C154 w_n7489_9836# a_1804_15931# 0.01614f
C155 w_n7489_9836# a_n7288_16809# 0.03158f
C156 m2_n74040_n58072# m3_n74040_n58072# 0.39453p
C157 a_5580_15247# a_n6059_11418# 0.66736f
C158 a_n7203_14433# a_n7289_16545# 0.28328f
C159 m5_n74040_n58072# m6_n74040_n58072# 0.25064p
C160 dw_n7489_9836# a_1804_15931# 5.15676f
C161 dw_n7489_9836# a_n7288_16809# 7.11994f
C162 a_3822_10479# a_3630_15211# 0.2774f
C163 m3_1900_17599# a_n6059_10861# 0.01692f
C164 a_n7202_17421# a_n6059_11418# 0.01101f
C165 w_3320_10081# a_3630_15211# 0.01456f
C166 a_527_16281# a_n7203_16545# 0.01946f
C167 a_5580_15247# a_3630_15211# 2.48993f
C168 a_n6059_11418# w_3320_16060# 0.0273f
C169 a_n7289_14961# a_n7203_14961# 0.01946f
C170 dw_n7489_9836# m3_1900_17599# 0.10215f
C171 a_n7203_16017# a_n7203_15753# 0.56632f
C172 a_n7289_14433# a_n7289_16545# 0.01035f
C173 a_3822_10479# w_8745_13831# 0.04005f
C174 m2_n73602_n57634# m1_n73602_n57634# 0.39413p
C175 a_3630_15211# w_3320_16060# 0.08623f
C176 a_n7289_16545# a_n7203_13669# 2.15576f
C177 w_1389_15644# a_n6059_11418# 0.01462f
C178 a_n7288_16809# a_n7288_17115# 0.0308f
C179 a_527_14697# a_n6059_10861# 0.0297f
C180 a_n7203_14697# a_n7289_16545# 0.27223f
C181 m3_1900_17599# a_1804_15931# 0.19321f
C182 a_n6059_11418# a_4707_16560# 1.8134f
C183 a_527_14697# a_n7289_16545# 0.01226f
C184 a_n7203_15225# a_n7203_14961# 0.56632f
C185 w_8745_13831# a_5580_15247# 0.01565f
C186 dw_n7489_9836# a_n7203_13669# 0.04526f
C187 a_527_15753# a_n7203_15753# 0.01946f
C188 a_n7202_17727# a_n7202_18033# 0.56632f
C189 a_n7203_16017# a_n7289_16545# 0.34937f
C190 a_n7202_18646# a_981_18638# 0.01155f
C191 w_1450_16710# a_n6059_10861# 0.01046f
C192 a_n7202_17727# a_n7288_17727# 0.02797f
C193 a_n7203_15489# a_n7289_15489# 0.01947f
C194 a_4707_16560# a_3630_15211# 2.47471f
C195 a_n7288_18340# dw_n7489_9836# 0.01497f
C196 a_n7288_16809# a_n7289_14433# 0.01845f
C197 m5_n73556_n57588# m4_n73602_n57634# 0.34892p
C198 a_527_15753# a_n6059_10861# 0.02893f
C199 a_n7288_16809# a_n7203_13669# 0.04028f
C200 dw_n7489_9836# w_1450_16710# 0.13974f
C201 a_n6059_11418# a_n6059_10861# 8.04164f
C202 m7_n74040_n58072# a_n74040_n58072# 0.19092p
C203 m6_n73460_n57492# a_n74040_n58072# 0.21787p
C204 m6_n74040_n58072# a_n74040_n58072# 0.21939p
C205 m5_n73556_n57588# a_n74040_n58072# 0.16053p
C206 m5_n74040_n58072# a_n74040_n58072# 0.16155p
C207 m4_n73602_n57634# a_n74040_n58072# 0.16966p
C208 m4_n74040_n58072# a_n74040_n58072# 0.17068p
C209 m3_1900_17599# a_n74040_n58072# 0.07285f
C210 m3_n73602_n57634# a_n74040_n58072# 0.1829p
C211 m3_n74040_n58072# a_n74040_n58072# 0.184p
C212 m2_n73602_n57634# a_n74040_n58072# 0.203p
C213 m2_n74040_n58072# a_n74040_n58072# 0.20422p
C214 m1_n73602_n57634# a_n74040_n58072# 0.43621p
C215 m1_n74040_n58072# a_n74040_n58072# 0.43781p
C216 a_n7059_10169# a_n74040_n58072# 18.9182f $ **FLOATING
C217 a_n7203_13669# a_n74040_n58072# 13.2663f
C218 a_527_13669# a_n74040_n58072# 0.57989f $ **FLOATING
C219 a_n7203_14433# a_n74040_n58072# 3.81224f
C220 a_n7203_14697# a_n74040_n58072# 3.80746f
C221 a_n7289_14433# a_n74040_n58072# 0.26883f $ **FLOATING
C222 a_3822_10479# a_n74040_n58072# 0.23654p $ **FLOATING
C223 a_527_14697# a_n74040_n58072# 0.25188f $ **FLOATING
C224 a_n7203_14961# a_n74040_n58072# 3.80233f
C225 a_n7203_15225# a_n74040_n58072# 3.79878f
C226 a_n7289_14961# a_n74040_n58072# 0.25151f $ **FLOATING
C227 a_n7203_15489# a_n74040_n58072# 3.79878f
C228 a_n7203_15753# a_n74040_n58072# 3.79878f
C229 a_n7289_15489# a_n74040_n58072# 0.25183f $ **FLOATING
C230 a_527_15753# a_n74040_n58072# 0.23297f $ **FLOATING
C231 a_n7203_16017# a_n74040_n58072# 3.79878f
C232 a_n7203_16281# a_n74040_n58072# 3.79878f
C233 a_n7289_16017# a_n74040_n58072# 0.25124f $ **FLOATING
C234 a_3630_15211# a_n74040_n58072# 6.36779f $ **FLOATING
C235 a_5580_15247# a_n74040_n58072# 51.4358f $ **FLOATING
C236 a_4707_16560# a_n74040_n58072# 1.69969f $ **FLOATING
C237 a_n6059_10861# a_n74040_n58072# 15.1337f $ **FLOATING
C238 a_1804_15931# a_n74040_n58072# 19.9354f $ **FLOATING
C239 a_n6059_11418# a_n74040_n58072# 9.66571f $ **FLOATING
C240 a_527_16281# a_n74040_n58072# 0.28604f $ **FLOATING
C241 a_n7203_16545# a_n74040_n58072# 3.79788f
C242 a_n7289_16545# a_n74040_n58072# 36.4829f $ **FLOATING
C243 a_n7202_16809# a_n74040_n58072# 4.50753f
C244 a_n7288_16809# a_n74040_n58072# 0.24344p $ **FLOATING
C245 a_528_16809# a_n74040_n58072# 0.34584f $ **FLOATING
C246 a_n7202_17115# a_n74040_n58072# 4.50921f
C247 a_n7202_17421# a_n74040_n58072# 4.50921f
C248 a_n7288_17115# a_n74040_n58072# 0.30345f $ **FLOATING
C249 a_528_17421# a_n74040_n58072# 0.34565f $ **FLOATING
C250 a_n7202_17727# a_n74040_n58072# 4.50921f
C251 a_n7202_18033# a_n74040_n58072# 4.51745f
C252 a_n7288_17727# a_n74040_n58072# 0.30438f $ **FLOATING
C253 a_528_18033# a_n74040_n58072# 0.36381f $ **FLOATING
C254 a_n7202_18340# a_n74040_n58072# 4.55105f
C255 a_981_18638# a_n74040_n58072# 1.17046f $ **FLOATING
C256 a_n7202_18646# a_n74040_n58072# 5.27974f
C257 a_n7288_18340# a_n74040_n58072# 0.3202f $ **FLOATING
C258 w_n7489_9836# a_n74040_n58072# 0.21456f
C259 w_3320_10081# a_n74040_n58072# 0.1031f
C260 w_8745_13831# a_n74040_n58072# 0.02418f
C261 w_3320_16060# a_n74040_n58072# 0.123f
C262 w_1450_16710# a_n74040_n58072# 0.03111f
C263 dw_n7489_9836# a_n74040_n58072# 0.52674p $ **FLOATING
.ends
