* Extracted by KLayout with SG13G2 LVS runset on : 10/07/2025 03:16

.SUBCKT ota_final
M$1 \$2 \$47 \$54 \$2 sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$5 \$2 \$47 \$47 \$2 sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$9 \$3 \$16 \$17 \$2 sg13_lv_nmos L=0.5u W=15u AS=3.4125p AD=3.4125p PS=20.57u
+ PD=20.57u
M$13 \$2 \$2 \$60 \$2 sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$14 \$60 \$67 \$53 \$2 sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p PS=6.76u
+ PD=6.76u
M$15 \$53 \$1 \$58 \$2 sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p PS=6.76u
+ PD=6.76u
M$16 \$58 \$2 \$2 \$2 sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$17 \$2 \$47 \$53 \$2 sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$25 \$54 \$46 \$56 \$3 sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p PS=19.32u
+ PD=19.32u
M$29 \$2 \$46 \$57 \$3 sg13_lv_pmos L=0.5u W=14u AS=3.185p AD=3.185p PS=19.32u
+ PD=19.32u
M$33 \$7 \$16 \$24 \$2 sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$35 \$2 \$2 \$7 \$2 sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$36 \$7 \$7 \$2 \$2 sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u PD=3.76u
M$37 \$2 \$7 \$17 \$2 sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u PD=3.76u
M$41 \$2 \$2 \$16 \$2 sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$42 \$16 \$17 \$I88 \$2 sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$45 \$2 \$2 \$I88 \$2 sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$46 \$I88 \$46 \$2 \$2 sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$49 \$2 \$2 \$I87 \$2 sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$50 \$I87 \$46 \$2 \$2 sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$53 \$2 \$2 \$46 \$2 sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$54 \$46 \$17 \$I87 \$2 sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$57 \$3 \$3 \$56 \$3 sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$58 \$56 \$56 \$3 \$3 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$59 \$3 \$56 \$57 \$3 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$61 \$3 \$56 \$24 \$3 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$71 \$3 \$3 \$46 \$3 sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$72 \$46 \$57 \$58 \$3 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$77 \$3 \$3 \$16 \$3 sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$78 \$16 \$57 \$60 \$3 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$83 \$3 \$3 \$60 \$3 sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p PS=19.32u
+ PD=19.32u
M$85 \$3 \$56 \$58 \$3 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$87 \$3 \$56 \$60 \$3 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
.ENDS ota_final
