.subckt analog_inverter VDD VSS
.ends
.end
