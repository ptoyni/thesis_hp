* Extracted by KLayout with SG13G2 LVS runset on : 21/08/2025 16:41

.SUBCKT foldedcascode_pmos AVDD AVSS IBIAS VOUT PLUS MINUS
M$1 AVSS AVSS \$45 AVSS sg13_lv_nmos L=2u W=1.33u AS=0.4522p AD=0.2527p
+ PS=3.34u PD=1.71u
M$2 \$45 \$22 \$33 AVSS sg13_lv_nmos L=2u W=1.33u AS=0.2527p AD=0.2527p
+ PS=1.71u PD=1.71u
M$3 \$33 AVSS AVSS AVSS sg13_lv_nmos L=2u W=5.33u AS=1.3127p AD=1.3127p
+ PS=8.77u PD=8.77u
M$4 AVSS AVSS \$36 AVSS sg13_lv_nmos L=2u W=1.33u AS=0.2527p AD=0.2527p
+ PS=1.71u PD=1.71u
M$5 \$36 \$22 VOUT AVSS sg13_lv_nmos L=2u W=1.33u AS=0.2527p AD=0.2527p
+ PS=1.71u PD=1.71u
M$6 VOUT AVSS AVSS AVSS sg13_lv_nmos L=2u W=1.33u AS=0.2527p AD=0.4522p
+ PS=1.71u PD=3.34u
C$7 VOUT AVSS cap_cmim w=25.82u l=25.82u A=666.6724p P=103.28u m=1
M$8 AVSS AVSS IBIAS AVSS sg13_lv_nmos L=2u W=4u AS=1.06p AD=1.06p PS=7.06u
+ PD=7.06u
M$9 IBIAS \$39 \$18 AVSS sg13_lv_nmos L=2u W=4u AS=0.76p AD=0.76p PS=4.76u
+ PD=4.76u
M$13 \$33 \$18 AVSS AVSS sg13_lv_nmos L=2u W=4u AS=0.76p AD=0.76p PS=4.76u
+ PD=4.76u
M$14 AVSS \$18 \$36 AVSS sg13_lv_nmos L=2u W=4u AS=0.76p AD=0.76p PS=4.76u
+ PD=4.76u
M$18 AVSS AVSS \$56 AVSS sg13_lv_nmos L=2u W=8u AS=2.12p AD=2.12p PS=13.06u
+ PD=13.06u
M$19 \$56 \$52 AVSS AVSS sg13_lv_nmos L=2u W=4u AS=0.76p AD=0.76p PS=4.38u
+ PD=4.38u
M$21 AVSS AVSS AVDD AVSS sg13_lv_nmos L=0.5u W=15u AS=3.975p AD=3.975p
+ PS=23.56u PD=23.56u
M$22 AVDD \$39 \$22 AVSS sg13_lv_nmos L=0.5u W=15u AS=2.85p AD=2.85p PS=15.76u
+ PD=15.76u
M$25 AVSS AVSS \$18 AVSS sg13_lv_nmos L=2u W=8u AS=2.12p AD=2.12p PS=13.06u
+ PD=13.06u
M$26 \$18 \$18 \$22 AVSS sg13_lv_nmos L=2u W=4u AS=0.76p AD=0.76p PS=4.38u
+ PD=4.38u
M$27 \$22 \$18 AVSS AVSS sg13_lv_nmos L=2u W=4u AS=0.76p AD=0.76p PS=4.38u
+ PD=4.38u
M$29 AVSS AVSS \$19 AVSS sg13_lv_nmos L=2u W=2u AS=0.68p AD=0.38p PS=4.68u
+ PD=2.38u
M$30 \$19 \$22 AVSS AVSS sg13_lv_nmos L=2u W=2u AS=0.38p AD=0.38p PS=2.38u
+ PD=2.38u
M$31 AVSS AVSS \$I231 AVSS sg13_lv_nmos L=2u W=2u AS=0.38p AD=0.68p PS=2.38u
+ PD=4.68u
M$32 AVDD AVDD \$56 AVDD sg13_lv_pmos L=5u W=14u AS=3.71p AD=3.71p PS=22.06u
+ PD=22.06u
M$33 \$56 \$56 AVDD AVDD sg13_lv_pmos L=5u W=28u AS=5.32p AD=5.32p PS=29.52u
+ PD=29.52u
M$38 AVDD AVDD AVDD AVDD sg13_lv_pmos L=5u W=16u AS=4.24p AD=4.24p PS=25.06u
+ PD=25.06u
M$39 AVDD \$56 \$77 AVDD sg13_lv_pmos L=5u W=32u AS=6.08p AD=6.08p PS=33.52u
+ PD=33.52u
M$44 AVDD AVDD \$77 AVDD sg13_lv_pmos L=2u W=20u AS=5.3p AD=5.3p PS=32.12u
+ PD=32.12u
M$45 \$77 PLUS \$33 AVDD sg13_lv_pmos L=2u W=20u AS=3.8p AD=3.8p PS=21.52u
+ PD=21.52u
M$47 \$77 MINUS \$36 AVDD sg13_lv_pmos L=2u W=20u AS=3.8p AD=3.8p PS=21.52u
+ PD=21.52u
M$56 \$34 \$34 \$19 AVDD sg13_lv_pmos L=2u W=4u AS=1.36p AD=0.76p PS=8.68u
+ PD=4.38u
M$57 \$19 \$19 \$I232 AVDD sg13_lv_pmos L=2u W=8u AS=1.52p AD=1.52p PS=8.76u
+ PD=8.76u
M$59 \$19 \$35 \$35 AVDD sg13_lv_pmos L=2u W=4u AS=0.76p AD=1.36p PS=4.38u
+ PD=8.68u
M$60 AVDD AVDD AVDD AVDD sg13_lv_pmos L=2u W=13u AS=3.445p AD=3.445p PS=20.56u
+ PD=20.56u
M$61 AVDD \$45 \$80 AVDD sg13_lv_pmos L=2u W=13u AS=2.47p AD=2.47p PS=13.76u
+ PD=13.76u
M$63 AVDD \$45 \$79 AVDD sg13_lv_pmos L=2u W=13u AS=2.47p AD=2.47p PS=13.76u
+ PD=13.76u
M$66 \$45 \$19 \$80 AVDD sg13_lv_pmos L=2u W=8u AS=2.72p AD=2.72p PS=16.68u
+ PD=16.68u
M$67 \$79 \$19 VOUT AVDD sg13_lv_pmos L=2u W=8u AS=2.72p AD=2.72p PS=16.68u
+ PD=16.68u
D$68 AVSS AVDD AVDD diodevdd_2kv m=1
D$69 AVSS AVDD AVSS diodevdd_2kv m=1
D$70 AVSS AVDD PLUS diodevdd_2kv m=1
D$71 AVSS AVDD VOUT diodevdd_2kv m=1
D$72 AVSS AVDD MINUS diodevdd_2kv m=1
D$73 AVSS AVDD IBIAS diodevdd_2kv m=1
D$74 AVDD AVSS MINUS diodevss_2kv m=1
D$75 AVDD AVSS IBIAS diodevss_2kv m=1
D$76 AVDD AVSS VOUT diodevss_2kv m=1
D$77 AVDD AVSS PLUS diodevss_2kv m=1
D$78 AVDD AVSS AVSS diodevss_2kv m=1
D$79 AVDD AVSS AVDD diodevss_2kv m=1
.ENDS foldedcascode_pmos
