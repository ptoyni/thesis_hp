* Extracted by KLayout with SG13G2 LVS runset on : 10/08/2025 02:57

.SUBCKT ota_final AVSS PLUS VOUT IBIAS MINUS
M$1 \$16463 VOUT \$18643 AVSS sg13_lv_nmos L=0.5u W=15u AS=3.4125p AD=3.4125p
+ PS=20.57u PD=20.57u
M$5 AVSS IBIAS IBIAS AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$9 AVSS IBIAS \$19588 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$13 AVSS IBIAS \$19587 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$17 AVSS AVSS \$19749 AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$18 \$19749 MINUS \$19587 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p
+ PS=6.76u PD=6.76u
M$19 \$19587 PLUS \$19750 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p
+ PS=6.76u PD=6.76u
M$20 \$19750 AVSS AVSS AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$25 \$19588 \$19073 \$19694 \$16463 sg13_lv_pmos L=2u W=14u AS=3.185p
+ AD=3.185p PS=19.32u PD=19.32u
M$29 AVSS \$19073 \$19695 \$16463 sg13_lv_pmos L=0.5u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
C$33 VOUT AVSS cap_cmim w=25.82u l=25.82u A=666.6724p P=103.28u m=1
M$34 \$18645 VOUT \$18646 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$36 AVSS AVSS \$18645 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$37 \$18645 \$18645 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$38 AVSS \$18645 \$18643 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$42 \$16463 \$16463 \$19694 \$16463 sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p
+ PS=11.56u PD=11.56u
M$43 \$19694 \$19694 \$16463 \$16463 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$44 \$16463 \$19694 \$19695 \$16463 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$46 \$16463 \$19694 \$18646 \$16463 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$56 AVSS AVSS VOUT AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$57 VOUT \$18643 \$I485994 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$60 AVSS AVSS \$I485993 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$61 \$I485993 \$19073 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$64 AVSS AVSS \$I485994 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$65 \$I485994 \$19073 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$68 AVSS AVSS \$19073 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$69 \$19073 \$18643 \$I485993 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$72 \$16463 \$16463 \$19073 \$16463 sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p
+ PS=11.56u PD=11.56u
M$73 \$19073 \$19695 \$19750 \$16463 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$78 \$16463 \$16463 VOUT \$16463 sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p
+ PS=11.56u PD=11.56u
M$79 VOUT \$19695 \$19749 \$16463 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$84 \$16463 \$16463 \$19749 \$16463 sg13_lv_pmos L=2u W=14u AS=3.185p
+ AD=3.185p PS=19.32u PD=19.32u
M$86 \$16463 \$19694 \$19750 \$16463 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$88 \$16463 \$19694 \$19749 \$16463 sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
.ENDS ota_final
