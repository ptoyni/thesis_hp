* Extracted by KLayout with SG13G2 LVS runset on : 25/05/2025 15:54

.SUBCKT analog_inverter VIN VOUT VDD VSS
M$1 VOUT VIN VSS \$5 sg13_lv_nmos L=0.52u W=1.3u AS=0.442p AD=0.442p PS=3.28u
+ PD=3.28u
M$2 VDD VIN VOUT \$I1 sg13_lv_pmos L=0.52u W=2.6u AS=0.884p AD=0.884p PS=5.88u
+ PD=5.88u
.ENDS analog_inverter
