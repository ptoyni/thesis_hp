* Extracted by KLayout with SG13G2 LVS runset on : 03/08/2025 21:18

.SUBCKT ota_final_decoup AVSS VOUT IBIAS MINUS PLUS AVDD
M$1 AVSS AVSS \$4 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$2 \$4 \$6 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u PD=3.76u
M$5 AVSS AVSS \$5 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$6 \$5 \$6 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u PD=3.76u
M$9 AVSS AVSS \$7 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$10 \$7 \$7 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$11 AVSS \$7 \$8 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$15 AVSS AVSS \$6 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$16 \$6 \$8 \$4 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u PD=3.76u
M$19 AVSS AVSS VOUT AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$20 VOUT \$8 \$5 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$23 AVDD VOUT \$8 AVSS sg13_lv_nmos L=0.5u W=15u AS=3.4125p AD=3.4125p
+ PS=20.57u PD=20.57u
M$27 AVSS IBIAS IBIAS AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$31 AVSS IBIAS \$19 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$35 AVSS IBIAS \$18 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$39 AVSS AVSS \$27 AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$40 \$27 MINUS \$18 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p PS=6.76u
+ PD=6.76u
M$41 \$18 PLUS \$21 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p PS=6.76u
+ PD=6.76u
M$42 \$21 AVSS AVSS AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$47 AVDD AVDD \$27 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p PS=19.32u
+ PD=19.32u
M$49 AVDD \$20 \$21 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$51 AVDD \$20 \$27 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$59 AVDD AVDD \$6 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$60 \$6 \$33 \$21 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$65 \$19 \$6 \$20 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p PS=19.32u
+ PD=19.32u
M$69 AVDD AVDD \$20 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$70 \$20 \$20 AVDD AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$71 AVDD \$20 \$33 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$73 AVDD \$20 \$34 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$83 AVSS \$6 \$33 AVDD sg13_lv_pmos L=0.5u W=14u AS=3.185p AD=3.185p PS=19.32u
+ PD=19.32u
M$87 AVDD AVDD VOUT AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$88 VOUT \$33 \$27 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$93 AVDD \$20 AVDD AVDD sg13_lv_pmos L=0.5u W=12u AS=2.73p AD=2.73p PS=16.82u
+ PD=16.82u
M$97 AVDD \$33 AVDD AVDD sg13_lv_pmos L=0.5u W=12u AS=2.73p AD=2.73p PS=16.82u
+ PD=16.82u
M$101 AVSS IBIAS AVSS AVSS sg13_lv_nmos L=1u W=8u AS=1.82p AD=1.82p PS=11.82u
+ PD=11.82u
M$105 AVSS \$8 AVSS AVSS sg13_lv_nmos L=1u W=8u AS=1.82p AD=1.82p PS=11.82u
+ PD=11.82u
C$109 VOUT AVSS cap_cmim w=25.82u l=25.82u A=666.6724p P=103.28u m=1
M$110 \$7 VOUT \$34 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
.ENDS ota_final_decoup
