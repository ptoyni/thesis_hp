* Extracted by KLayout with SG13G2 LVS runset on : 22/08/2025 15:02

.SUBCKT ota_final AVDD IBIAS VOUT MINUS PLUS AVSS
XM1 AVSS AVSS \$20 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
XM2 \$20 \$22 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
XM5 AVSS AVSS \$21 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
XM6 \$21 \$22 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
XM9 AVSS AVSS \$23 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
XM10 \$23 \$23 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
XM11 AVSS \$23 \$25 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
XM15 AVSS AVSS \$22 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
XM16 \$22 \$25 \$20 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
XM19 AVSS AVSS VOUT AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
XM20 VOUT \$25 \$21 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
XM23 AVDD VOUT \$25 AVSS sg13_lv_nmos L=0.5u W=15u AS=3.4125p AD=3.4125p
+ PS=20.57u PD=20.57u
XM27 AVSS IBIAS IBIAS AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
XM31 AVSS IBIAS \$36 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
XM35 AVSS IBIAS \$35 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
XM39 AVSS AVSS \$44 AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
XM40 \$44 MINUS \$35 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p PS=6.76u
+ PD=6.76u
XM41 \$35 PLUS \$38 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p PS=6.76u
+ PD=6.76u
XM42 \$38 AVSS AVSS AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
XM47 AVDD AVDD \$44 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p PS=19.32u
+ PD=19.32u
XM49 AVDD \$37 \$38 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
XM51 AVDD \$37 \$44 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
XM59 AVDD AVDD \$22 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
XM60 \$22 \$51 \$38 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
XM65 \$36 \$22 \$37 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p PS=19.32u
+ PD=19.32u
XM69 AVDD AVDD \$37 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
XM70 \$37 \$37 AVDD AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
XM71 AVDD \$37 \$51 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
XM73 AVDD \$37 \$52 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
XM83 AVSS \$22 \$51 AVDD sg13_lv_pmos L=0.5u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
XM87 AVDD AVDD VOUT AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
XM88 VOUT \$51 \$44 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
XM93 AVDD \$37 AVDD AVDD sg13_lv_pmos L=0.5u W=12u AS=2.73p AD=2.73p PS=16.82u
+ PD=16.82u
XM97 AVDD \$51 AVDD AVDD sg13_lv_pmos L=0.5u W=12u AS=2.73p AD=2.73p PS=16.82u
+ PD=16.82u
XM101 AVSS IBIAS AVSS AVSS sg13_lv_nmos L=1u W=8u AS=1.82p AD=1.82p PS=11.82u
+ PD=11.82u
XM105 AVSS \$25 AVSS AVSS sg13_lv_nmos L=1u W=8u AS=1.82p AD=1.82p PS=11.82u
+ PD=11.82u
XC115 VOUT AVSS cap_cmim w=25.82u l=25.82u A=666.6724p P=103.28u m=1
XM116 \$23 VOUT \$52 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
.ENDS FMD_QNC_ota_decoup
