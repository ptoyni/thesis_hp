* Extracted by KLayout with SG13G2 LVS runset on : 05/07/2025 18:36

.SUBCKT foldedcascode_nmos_withdummies AVSS D_ENA VOUT IBIAS AVDD PLUS MINUS
M$1 AVSS \$3 \$2 AVSS sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$2 AVSS AVSS \$65 AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$3 \$65 PLUS \$60 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p PS=6.76u
+ PD=6.76u
M$4 \$60 MINUS \$70 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p PS=6.76u
+ PD=6.76u
M$5 \$70 AVSS AVSS AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$10 IBIAS \$51 \$52 AVSS sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$11 AVSS VOUT \$20 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$13 AVDD VOUT \$12 AVSS sg13_lv_nmos L=0.5u W=15u AS=3.4125p AD=3.4125p
+ PS=20.57u PD=20.57u
M$17 AVSS \$68 \$67 AVDD sg13_lv_pmos L=0.5u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
M$21 \$61 \$68 \$66 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p PS=19.32u
+ PD=19.32u
M$25 AVSS \$3 \$51 AVSS sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$26 AVSS D_ENA \$3 AVSS sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$27 AVDD \$3 \$51 AVDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$28 AVDD D_ENA \$3 AVDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$29 AVSS \$52 IBIAS AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$33 AVSS \$52 \$60 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$37 AVSS \$52 \$53 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$41 AVSS AVSS \$I49 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$42 \$I49 \$I49 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$43 AVSS \$I49 \$12 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$47 AVSS AVSS VOUT AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$48 VOUT \$12 \$I52 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$51 AVSS AVSS \$I50 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$52 \$I50 \$2 \$I51 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$55 AVSS AVSS \$I52 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$56 \$I52 \$2 \$I53 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$59 AVSS AVSS \$2 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$60 \$2 \$12 \$I50 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p PS=3.76u
+ PD=3.76u
M$63 AVDD AVDD \$66 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$64 \$66 \$66 AVDD AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$65 AVDD \$66 \$67 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$67 AVDD \$66 \$20 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$77 AVDD AVDD \$2 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$78 \$2 \$67 \$70 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$83 AVDD AVDD VOUT AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$84 VOUT \$67 \$65 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$89 AVDD AVDD \$65 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p PS=19.32u
+ PD=19.32u
M$91 AVDD \$66 \$70 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$93 AVDD \$66 \$65 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p PS=15.52u
+ PD=15.52u
M$101 AVDD \$67 AVDD AVDD sg13_lv_pmos L=1u W=64u AS=14.56p AD=14.56p PS=83.64u
+ PD=83.64u
M$109 AVSS \$12 AVSS AVSS sg13_lv_nmos L=1u W=32u AS=7.28p AD=7.28p PS=41.82u
+ PD=41.82u
M$113 AVSS \$60 AVSS AVSS sg13_lv_nmos L=1u W=32u AS=7.28p AD=7.28p PS=41.82u
+ PD=41.82u
.ENDS foldedcascode_nmos_withdummies
