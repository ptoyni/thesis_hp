* Extracted by KLayout with SG13G2 LVS runset on : 11/07/2025 16:52

.SUBCKT ota_final AVSS PLUS IBIAS AVDD VOUT MINUS
M$1 AVDD VOUT \$18329 AVSS sg13_lv_nmos L=0.5u W=15u AS=3.4125p AD=3.4125p
+ PS=20.57u PD=20.57u
M$5 AVSS IBIAS IBIAS AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$9 AVSS IBIAS \$19325 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$13 AVSS IBIAS \$19324 AVSS sg13_lv_nmos L=5u W=8.5u AS=1.93375p AD=1.93375p
+ PS=12.445u PD=12.445u
M$17 AVSS AVSS \$19436 AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$18 \$19436 MINUS \$19324 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p
+ PS=6.76u PD=6.76u
M$19 \$19324 PLUS \$19652 AVSS sg13_lv_nmos L=1u W=6u AS=1.14p AD=1.14p
+ PS=6.76u PD=6.76u
M$20 \$19652 AVSS AVSS AVSS sg13_lv_nmos L=1u W=6u AS=1.59p AD=1.59p PS=10.06u
+ PD=10.06u
M$25 \$19325 \$18745 \$19326 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
M$29 AVSS \$18745 \$19328 AVDD sg13_lv_pmos L=0.5u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
M$33 \$18331 VOUT \$18467 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$35 AVSS AVSS \$18331 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$36 \$18331 \$18331 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$37 AVSS \$18331 \$18329 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$41 AVSS AVSS VOUT AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$42 VOUT \$18329 \$I498845 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$45 AVSS AVSS \$I498844 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$46 \$I498844 \$18745 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$49 AVSS AVSS \$I498845 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p
+ PS=5.56u PD=5.56u
M$50 \$I498845 \$18745 AVSS AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$53 AVSS AVSS \$18745 AVSS sg13_lv_nmos L=2u W=3u AS=0.795p AD=0.795p PS=5.56u
+ PD=5.56u
M$54 \$18745 \$18329 \$I498844 AVSS sg13_lv_nmos L=2u W=3u AS=0.57p AD=0.57p
+ PS=3.76u PD=3.76u
M$57 AVDD AVDD \$19326 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p
+ PS=11.56u PD=11.56u
M$58 \$19326 \$19326 AVDD AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$59 AVDD \$19326 \$19328 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$61 AVDD \$19326 \$18467 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$71 AVDD AVDD \$18745 AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p
+ PS=11.56u PD=11.56u
M$72 \$18745 \$19328 \$19652 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$77 AVDD AVDD VOUT AVDD sg13_lv_pmos L=2u W=7u AS=1.855p AD=1.855p PS=11.56u
+ PD=11.56u
M$78 VOUT \$19328 \$19436 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$83 AVDD AVDD \$19436 AVDD sg13_lv_pmos L=2u W=14u AS=3.185p AD=3.185p
+ PS=19.32u PD=19.32u
M$85 AVDD \$19326 \$19652 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
M$87 AVDD \$19326 \$19436 AVDD sg13_lv_pmos L=2u W=14u AS=2.66p AD=2.66p
+ PS=15.52u PD=15.52u
.ENDS ota_final
