.SUBCKT analog_inverter VIN VOUT VDD VSS
*.ipin VIN
*.iopin VDD
*.iopin VSS
*.opin VOUT
MN1 VOUT VIN VSS VSS sg13_lv_nmos w=1.3u l=0.52u ng=1 m=1
MP1 VOUT VIN VDD VDD sg13_lv_pmos w=2.6u l=0.52u ng=1 m=1
.ENDS