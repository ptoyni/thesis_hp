** sch_path: /foss/designs/thesis/workspace/thesis_hp/Designs/Analog_Inverter/Schematics/Analog_Inverter.sch
**.subckt Analog_Inverter vdd vin vout vss
*.ipin vin
*.iopin vdd
*.iopin vss
*.opin vout
XM1 vout vin vdd vdd sg13_lv_pmos w=2u l=0.15u ng=1 m=1
XM2 vout vin vss vss sg13_lv_nmos w=1u l=0.15u ng=1 m=1
**.ends
.end
