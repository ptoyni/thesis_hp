* Extracted by KLayout with SG13G2 LVS runset on : 29/06/2025 21:42

.SUBCKT enable_pins vss D_ENA AVDD
M$1 \$4 \$3 vss vss sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$2 \$4 \$3 AVDD AVDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$3 \$3 D_ENA vss vss sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$4 \$3 D_ENA AVDD AVDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
.ENDS enable_pins
