** sch_path: /foss/designs/thesis/workspace/thesis_hp/designs/analog_inverter/1_schematics/Analog_Inverter.sch
.subckt Analog_Inverter vdd vin vout vss
*.PININFO vin:I vdd:B vss:B vout:O
M1 vout vin vdd vdd sg13_lv_pmos w=2.6u l=0.52u ng=1 m=1
M2 vout vin vss vss sg13_lv_nmos w=1.3u l=0.52u ng=1 m=1
.ends
